module Arbiter(
  input          io_in_0_valid,
  input  [34:0]  io_in_0_bits_waddr,
  input  [4:0]   io_in_0_bits_entryid,
  input  [13:0]  io_in_0_bits_awid,
  input  [255:0] io_in_0_bits_data,
  input  [31:0]  io_in_0_bits_mask,
  input  [2:0]   io_in_0_bits_size,
  input  [7:0]   io_in_0_bits_len,
  input          io_in_1_valid,
  input  [34:0]  io_in_1_bits_waddr,
  input  [4:0]   io_in_1_bits_entryid,
  input  [13:0]  io_in_1_bits_awid,
  input  [255:0] io_in_1_bits_data,
  input  [31:0]  io_in_1_bits_mask,
  input  [2:0]   io_in_1_bits_size,
  input  [7:0]   io_in_1_bits_len,
  input          io_in_2_valid,
  input  [34:0]  io_in_2_bits_waddr,
  input  [4:0]   io_in_2_bits_entryid,
  input  [13:0]  io_in_2_bits_awid,
  input  [255:0] io_in_2_bits_data,
  input  [31:0]  io_in_2_bits_mask,
  input  [2:0]   io_in_2_bits_size,
  input  [7:0]   io_in_2_bits_len,
  input          io_in_3_valid,
  input  [34:0]  io_in_3_bits_waddr,
  input  [4:0]   io_in_3_bits_entryid,
  input  [13:0]  io_in_3_bits_awid,
  input  [255:0] io_in_3_bits_data,
  input  [31:0]  io_in_3_bits_mask,
  input  [2:0]   io_in_3_bits_size,
  input  [7:0]   io_in_3_bits_len,
  input          io_in_4_valid,
  input  [34:0]  io_in_4_bits_waddr,
  input  [4:0]   io_in_4_bits_entryid,
  input  [13:0]  io_in_4_bits_awid,
  input  [255:0] io_in_4_bits_data,
  input  [31:0]  io_in_4_bits_mask,
  input  [2:0]   io_in_4_bits_size,
  input  [7:0]   io_in_4_bits_len,
  input          io_in_5_valid,
  input  [34:0]  io_in_5_bits_waddr,
  input  [4:0]   io_in_5_bits_entryid,
  input  [13:0]  io_in_5_bits_awid,
  input  [255:0] io_in_5_bits_data,
  input  [31:0]  io_in_5_bits_mask,
  input  [2:0]   io_in_5_bits_size,
  input  [7:0]   io_in_5_bits_len,
  input          io_in_6_valid,
  input  [34:0]  io_in_6_bits_waddr,
  input  [4:0]   io_in_6_bits_entryid,
  input  [13:0]  io_in_6_bits_awid,
  input  [255:0] io_in_6_bits_data,
  input  [31:0]  io_in_6_bits_mask,
  input  [2:0]   io_in_6_bits_size,
  input  [7:0]   io_in_6_bits_len,
  input          io_in_7_valid,
  input  [34:0]  io_in_7_bits_waddr,
  input  [4:0]   io_in_7_bits_entryid,
  input  [13:0]  io_in_7_bits_awid,
  input  [255:0] io_in_7_bits_data,
  input  [31:0]  io_in_7_bits_mask,
  input  [2:0]   io_in_7_bits_size,
  input  [7:0]   io_in_7_bits_len,
  input          io_in_8_valid,
  input  [34:0]  io_in_8_bits_waddr,
  input  [4:0]   io_in_8_bits_entryid,
  input  [13:0]  io_in_8_bits_awid,
  input  [255:0] io_in_8_bits_data,
  input  [31:0]  io_in_8_bits_mask,
  input  [2:0]   io_in_8_bits_size,
  input  [7:0]   io_in_8_bits_len,
  input          io_in_9_valid,
  input  [34:0]  io_in_9_bits_waddr,
  input  [4:0]   io_in_9_bits_entryid,
  input  [13:0]  io_in_9_bits_awid,
  input  [255:0] io_in_9_bits_data,
  input  [31:0]  io_in_9_bits_mask,
  input  [2:0]   io_in_9_bits_size,
  input  [7:0]   io_in_9_bits_len,
  input          io_in_10_valid,
  input  [34:0]  io_in_10_bits_waddr,
  input  [4:0]   io_in_10_bits_entryid,
  input  [13:0]  io_in_10_bits_awid,
  input  [255:0] io_in_10_bits_data,
  input  [31:0]  io_in_10_bits_mask,
  input  [2:0]   io_in_10_bits_size,
  input  [7:0]   io_in_10_bits_len,
  input          io_in_11_valid,
  input  [34:0]  io_in_11_bits_waddr,
  input  [4:0]   io_in_11_bits_entryid,
  input  [13:0]  io_in_11_bits_awid,
  input  [255:0] io_in_11_bits_data,
  input  [31:0]  io_in_11_bits_mask,
  input  [2:0]   io_in_11_bits_size,
  input  [7:0]   io_in_11_bits_len,
  input          io_in_12_valid,
  input  [34:0]  io_in_12_bits_waddr,
  input  [4:0]   io_in_12_bits_entryid,
  input  [13:0]  io_in_12_bits_awid,
  input  [255:0] io_in_12_bits_data,
  input  [31:0]  io_in_12_bits_mask,
  input  [2:0]   io_in_12_bits_size,
  input  [7:0]   io_in_12_bits_len,
  input          io_in_13_valid,
  input  [34:0]  io_in_13_bits_waddr,
  input  [4:0]   io_in_13_bits_entryid,
  input  [13:0]  io_in_13_bits_awid,
  input  [255:0] io_in_13_bits_data,
  input  [31:0]  io_in_13_bits_mask,
  input  [2:0]   io_in_13_bits_size,
  input  [7:0]   io_in_13_bits_len,
  input          io_in_14_valid,
  input  [34:0]  io_in_14_bits_waddr,
  input  [4:0]   io_in_14_bits_entryid,
  input  [13:0]  io_in_14_bits_awid,
  input  [255:0] io_in_14_bits_data,
  input  [31:0]  io_in_14_bits_mask,
  input  [2:0]   io_in_14_bits_size,
  input  [7:0]   io_in_14_bits_len,
  input          io_in_15_valid,
  input  [34:0]  io_in_15_bits_waddr,
  input  [4:0]   io_in_15_bits_entryid,
  input  [13:0]  io_in_15_bits_awid,
  input  [255:0] io_in_15_bits_data,
  input  [31:0]  io_in_15_bits_mask,
  input  [2:0]   io_in_15_bits_size,
  input  [7:0]   io_in_15_bits_len,
  input          io_in_16_valid,
  input  [34:0]  io_in_16_bits_waddr,
  input  [4:0]   io_in_16_bits_entryid,
  input  [13:0]  io_in_16_bits_awid,
  input  [255:0] io_in_16_bits_data,
  input  [31:0]  io_in_16_bits_mask,
  input  [2:0]   io_in_16_bits_size,
  input  [7:0]   io_in_16_bits_len,
  input          io_in_17_valid,
  input  [34:0]  io_in_17_bits_waddr,
  input  [4:0]   io_in_17_bits_entryid,
  input  [13:0]  io_in_17_bits_awid,
  input  [255:0] io_in_17_bits_data,
  input  [31:0]  io_in_17_bits_mask,
  input  [2:0]   io_in_17_bits_size,
  input  [7:0]   io_in_17_bits_len,
  input          io_in_18_valid,
  input  [34:0]  io_in_18_bits_waddr,
  input  [4:0]   io_in_18_bits_entryid,
  input  [13:0]  io_in_18_bits_awid,
  input  [255:0] io_in_18_bits_data,
  input  [31:0]  io_in_18_bits_mask,
  input  [2:0]   io_in_18_bits_size,
  input  [7:0]   io_in_18_bits_len,
  input          io_in_19_valid,
  input  [34:0]  io_in_19_bits_waddr,
  input  [4:0]   io_in_19_bits_entryid,
  input  [13:0]  io_in_19_bits_awid,
  input  [255:0] io_in_19_bits_data,
  input  [31:0]  io_in_19_bits_mask,
  input  [2:0]   io_in_19_bits_size,
  input  [7:0]   io_in_19_bits_len,
  input          io_in_20_valid,
  input  [34:0]  io_in_20_bits_waddr,
  input  [4:0]   io_in_20_bits_entryid,
  input  [13:0]  io_in_20_bits_awid,
  input  [255:0] io_in_20_bits_data,
  input  [31:0]  io_in_20_bits_mask,
  input  [2:0]   io_in_20_bits_size,
  input  [7:0]   io_in_20_bits_len,
  input          io_in_21_valid,
  input  [34:0]  io_in_21_bits_waddr,
  input  [4:0]   io_in_21_bits_entryid,
  input  [13:0]  io_in_21_bits_awid,
  input  [255:0] io_in_21_bits_data,
  input  [31:0]  io_in_21_bits_mask,
  input  [2:0]   io_in_21_bits_size,
  input  [7:0]   io_in_21_bits_len,
  input          io_in_22_valid,
  input  [34:0]  io_in_22_bits_waddr,
  input  [4:0]   io_in_22_bits_entryid,
  input  [13:0]  io_in_22_bits_awid,
  input  [255:0] io_in_22_bits_data,
  input  [31:0]  io_in_22_bits_mask,
  input  [2:0]   io_in_22_bits_size,
  input  [7:0]   io_in_22_bits_len,
  input          io_in_23_valid,
  input  [34:0]  io_in_23_bits_waddr,
  input  [4:0]   io_in_23_bits_entryid,
  input  [13:0]  io_in_23_bits_awid,
  input  [255:0] io_in_23_bits_data,
  input  [31:0]  io_in_23_bits_mask,
  input  [2:0]   io_in_23_bits_size,
  input  [7:0]   io_in_23_bits_len,
  input          io_in_24_valid,
  input  [34:0]  io_in_24_bits_waddr,
  input  [4:0]   io_in_24_bits_entryid,
  input  [13:0]  io_in_24_bits_awid,
  input  [255:0] io_in_24_bits_data,
  input  [31:0]  io_in_24_bits_mask,
  input  [2:0]   io_in_24_bits_size,
  input  [7:0]   io_in_24_bits_len,
  input          io_in_25_valid,
  input  [34:0]  io_in_25_bits_waddr,
  input  [4:0]   io_in_25_bits_entryid,
  input  [13:0]  io_in_25_bits_awid,
  input  [255:0] io_in_25_bits_data,
  input  [31:0]  io_in_25_bits_mask,
  input  [2:0]   io_in_25_bits_size,
  input  [7:0]   io_in_25_bits_len,
  input          io_in_26_valid,
  input  [34:0]  io_in_26_bits_waddr,
  input  [4:0]   io_in_26_bits_entryid,
  input  [13:0]  io_in_26_bits_awid,
  input  [255:0] io_in_26_bits_data,
  input  [31:0]  io_in_26_bits_mask,
  input  [2:0]   io_in_26_bits_size,
  input  [7:0]   io_in_26_bits_len,
  input          io_in_27_valid,
  input  [34:0]  io_in_27_bits_waddr,
  input  [4:0]   io_in_27_bits_entryid,
  input  [13:0]  io_in_27_bits_awid,
  input  [255:0] io_in_27_bits_data,
  input  [31:0]  io_in_27_bits_mask,
  input  [2:0]   io_in_27_bits_size,
  input  [7:0]   io_in_27_bits_len,
  input          io_in_28_valid,
  input  [34:0]  io_in_28_bits_waddr,
  input  [4:0]   io_in_28_bits_entryid,
  input  [13:0]  io_in_28_bits_awid,
  input  [255:0] io_in_28_bits_data,
  input  [31:0]  io_in_28_bits_mask,
  input  [2:0]   io_in_28_bits_size,
  input  [7:0]   io_in_28_bits_len,
  input          io_in_29_valid,
  input  [34:0]  io_in_29_bits_waddr,
  input  [4:0]   io_in_29_bits_entryid,
  input  [13:0]  io_in_29_bits_awid,
  input  [255:0] io_in_29_bits_data,
  input  [31:0]  io_in_29_bits_mask,
  input  [2:0]   io_in_29_bits_size,
  input  [7:0]   io_in_29_bits_len,
  input          io_in_30_valid,
  input  [34:0]  io_in_30_bits_waddr,
  input  [4:0]   io_in_30_bits_entryid,
  input  [13:0]  io_in_30_bits_awid,
  input  [255:0] io_in_30_bits_data,
  input  [31:0]  io_in_30_bits_mask,
  input  [2:0]   io_in_30_bits_size,
  input  [7:0]   io_in_30_bits_len,
  input          io_in_31_valid,
  input  [34:0]  io_in_31_bits_waddr,
  input  [4:0]   io_in_31_bits_entryid,
  input  [13:0]  io_in_31_bits_awid,
  input  [255:0] io_in_31_bits_data,
  input  [31:0]  io_in_31_bits_mask,
  input  [2:0]   io_in_31_bits_size,
  input  [7:0]   io_in_31_bits_len,
  output         io_out_valid,
  output [34:0]  io_out_bits_waddr,
  output [4:0]   io_out_bits_entryid,
  output [13:0]  io_out_bits_awid,
  output [255:0] io_out_bits_data,
  output [31:0]  io_out_bits_mask,
  output [2:0]   io_out_bits_size,
  output [7:0]   io_out_bits_len
);
  wire [7:0] _GEN_1 = io_in_30_valid ? io_in_30_bits_len : io_in_31_bits_len; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [2:0] _GEN_2 = io_in_30_valid ? io_in_30_bits_size : io_in_31_bits_size; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [31:0] _GEN_4 = io_in_30_valid ? io_in_30_bits_mask : io_in_31_bits_mask; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [255:0] _GEN_5 = io_in_30_valid ? io_in_30_bits_data : io_in_31_bits_data; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [13:0] _GEN_12 = io_in_30_valid ? io_in_30_bits_awid : io_in_31_bits_awid; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [4:0] _GEN_13 = io_in_30_valid ? io_in_30_bits_entryid : io_in_31_bits_entryid; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [34:0] _GEN_16 = io_in_30_valid ? io_in_30_bits_waddr : io_in_31_bits_waddr; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [7:0] _GEN_20 = io_in_29_valid ? io_in_29_bits_len : _GEN_1; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_21 = io_in_29_valid ? io_in_29_bits_size : _GEN_2; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_23 = io_in_29_valid ? io_in_29_bits_mask : _GEN_4; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_24 = io_in_29_valid ? io_in_29_bits_data : _GEN_5; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_31 = io_in_29_valid ? io_in_29_bits_awid : _GEN_12; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_32 = io_in_29_valid ? io_in_29_bits_entryid : _GEN_13; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_35 = io_in_29_valid ? io_in_29_bits_waddr : _GEN_16; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_39 = io_in_28_valid ? io_in_28_bits_len : _GEN_20; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_40 = io_in_28_valid ? io_in_28_bits_size : _GEN_21; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_42 = io_in_28_valid ? io_in_28_bits_mask : _GEN_23; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_43 = io_in_28_valid ? io_in_28_bits_data : _GEN_24; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_50 = io_in_28_valid ? io_in_28_bits_awid : _GEN_31; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_51 = io_in_28_valid ? io_in_28_bits_entryid : _GEN_32; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_54 = io_in_28_valid ? io_in_28_bits_waddr : _GEN_35; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_58 = io_in_27_valid ? io_in_27_bits_len : _GEN_39; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_59 = io_in_27_valid ? io_in_27_bits_size : _GEN_40; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_61 = io_in_27_valid ? io_in_27_bits_mask : _GEN_42; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_62 = io_in_27_valid ? io_in_27_bits_data : _GEN_43; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_69 = io_in_27_valid ? io_in_27_bits_awid : _GEN_50; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_70 = io_in_27_valid ? io_in_27_bits_entryid : _GEN_51; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_73 = io_in_27_valid ? io_in_27_bits_waddr : _GEN_54; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_77 = io_in_26_valid ? io_in_26_bits_len : _GEN_58; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_78 = io_in_26_valid ? io_in_26_bits_size : _GEN_59; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_80 = io_in_26_valid ? io_in_26_bits_mask : _GEN_61; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_81 = io_in_26_valid ? io_in_26_bits_data : _GEN_62; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_88 = io_in_26_valid ? io_in_26_bits_awid : _GEN_69; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_89 = io_in_26_valid ? io_in_26_bits_entryid : _GEN_70; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_92 = io_in_26_valid ? io_in_26_bits_waddr : _GEN_73; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_96 = io_in_25_valid ? io_in_25_bits_len : _GEN_77; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_97 = io_in_25_valid ? io_in_25_bits_size : _GEN_78; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_99 = io_in_25_valid ? io_in_25_bits_mask : _GEN_80; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_100 = io_in_25_valid ? io_in_25_bits_data : _GEN_81; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_107 = io_in_25_valid ? io_in_25_bits_awid : _GEN_88; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_108 = io_in_25_valid ? io_in_25_bits_entryid : _GEN_89; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_111 = io_in_25_valid ? io_in_25_bits_waddr : _GEN_92; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_115 = io_in_24_valid ? io_in_24_bits_len : _GEN_96; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_116 = io_in_24_valid ? io_in_24_bits_size : _GEN_97; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_118 = io_in_24_valid ? io_in_24_bits_mask : _GEN_99; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_119 = io_in_24_valid ? io_in_24_bits_data : _GEN_100; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_126 = io_in_24_valid ? io_in_24_bits_awid : _GEN_107; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_127 = io_in_24_valid ? io_in_24_bits_entryid : _GEN_108; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_130 = io_in_24_valid ? io_in_24_bits_waddr : _GEN_111; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_134 = io_in_23_valid ? io_in_23_bits_len : _GEN_115; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_135 = io_in_23_valid ? io_in_23_bits_size : _GEN_116; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_137 = io_in_23_valid ? io_in_23_bits_mask : _GEN_118; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_138 = io_in_23_valid ? io_in_23_bits_data : _GEN_119; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_145 = io_in_23_valid ? io_in_23_bits_awid : _GEN_126; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_146 = io_in_23_valid ? io_in_23_bits_entryid : _GEN_127; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_149 = io_in_23_valid ? io_in_23_bits_waddr : _GEN_130; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_153 = io_in_22_valid ? io_in_22_bits_len : _GEN_134; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_154 = io_in_22_valid ? io_in_22_bits_size : _GEN_135; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_156 = io_in_22_valid ? io_in_22_bits_mask : _GEN_137; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_157 = io_in_22_valid ? io_in_22_bits_data : _GEN_138; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_164 = io_in_22_valid ? io_in_22_bits_awid : _GEN_145; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_165 = io_in_22_valid ? io_in_22_bits_entryid : _GEN_146; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_168 = io_in_22_valid ? io_in_22_bits_waddr : _GEN_149; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_172 = io_in_21_valid ? io_in_21_bits_len : _GEN_153; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_173 = io_in_21_valid ? io_in_21_bits_size : _GEN_154; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_175 = io_in_21_valid ? io_in_21_bits_mask : _GEN_156; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_176 = io_in_21_valid ? io_in_21_bits_data : _GEN_157; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_183 = io_in_21_valid ? io_in_21_bits_awid : _GEN_164; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_184 = io_in_21_valid ? io_in_21_bits_entryid : _GEN_165; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_187 = io_in_21_valid ? io_in_21_bits_waddr : _GEN_168; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_191 = io_in_20_valid ? io_in_20_bits_len : _GEN_172; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_192 = io_in_20_valid ? io_in_20_bits_size : _GEN_173; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_194 = io_in_20_valid ? io_in_20_bits_mask : _GEN_175; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_195 = io_in_20_valid ? io_in_20_bits_data : _GEN_176; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_202 = io_in_20_valid ? io_in_20_bits_awid : _GEN_183; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_203 = io_in_20_valid ? io_in_20_bits_entryid : _GEN_184; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_206 = io_in_20_valid ? io_in_20_bits_waddr : _GEN_187; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_210 = io_in_19_valid ? io_in_19_bits_len : _GEN_191; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_211 = io_in_19_valid ? io_in_19_bits_size : _GEN_192; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_213 = io_in_19_valid ? io_in_19_bits_mask : _GEN_194; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_214 = io_in_19_valid ? io_in_19_bits_data : _GEN_195; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_221 = io_in_19_valid ? io_in_19_bits_awid : _GEN_202; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_222 = io_in_19_valid ? io_in_19_bits_entryid : _GEN_203; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_225 = io_in_19_valid ? io_in_19_bits_waddr : _GEN_206; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_229 = io_in_18_valid ? io_in_18_bits_len : _GEN_210; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_230 = io_in_18_valid ? io_in_18_bits_size : _GEN_211; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_232 = io_in_18_valid ? io_in_18_bits_mask : _GEN_213; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_233 = io_in_18_valid ? io_in_18_bits_data : _GEN_214; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_240 = io_in_18_valid ? io_in_18_bits_awid : _GEN_221; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_241 = io_in_18_valid ? io_in_18_bits_entryid : _GEN_222; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_244 = io_in_18_valid ? io_in_18_bits_waddr : _GEN_225; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_248 = io_in_17_valid ? io_in_17_bits_len : _GEN_229; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_249 = io_in_17_valid ? io_in_17_bits_size : _GEN_230; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_251 = io_in_17_valid ? io_in_17_bits_mask : _GEN_232; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_252 = io_in_17_valid ? io_in_17_bits_data : _GEN_233; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_259 = io_in_17_valid ? io_in_17_bits_awid : _GEN_240; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_260 = io_in_17_valid ? io_in_17_bits_entryid : _GEN_241; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_263 = io_in_17_valid ? io_in_17_bits_waddr : _GEN_244; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_267 = io_in_16_valid ? io_in_16_bits_len : _GEN_248; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_268 = io_in_16_valid ? io_in_16_bits_size : _GEN_249; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_270 = io_in_16_valid ? io_in_16_bits_mask : _GEN_251; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_271 = io_in_16_valid ? io_in_16_bits_data : _GEN_252; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_278 = io_in_16_valid ? io_in_16_bits_awid : _GEN_259; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_279 = io_in_16_valid ? io_in_16_bits_entryid : _GEN_260; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_282 = io_in_16_valid ? io_in_16_bits_waddr : _GEN_263; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_286 = io_in_15_valid ? io_in_15_bits_len : _GEN_267; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_287 = io_in_15_valid ? io_in_15_bits_size : _GEN_268; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_289 = io_in_15_valid ? io_in_15_bits_mask : _GEN_270; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_290 = io_in_15_valid ? io_in_15_bits_data : _GEN_271; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_297 = io_in_15_valid ? io_in_15_bits_awid : _GEN_278; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_298 = io_in_15_valid ? io_in_15_bits_entryid : _GEN_279; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_301 = io_in_15_valid ? io_in_15_bits_waddr : _GEN_282; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_305 = io_in_14_valid ? io_in_14_bits_len : _GEN_286; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_306 = io_in_14_valid ? io_in_14_bits_size : _GEN_287; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_308 = io_in_14_valid ? io_in_14_bits_mask : _GEN_289; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_309 = io_in_14_valid ? io_in_14_bits_data : _GEN_290; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_316 = io_in_14_valid ? io_in_14_bits_awid : _GEN_297; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_317 = io_in_14_valid ? io_in_14_bits_entryid : _GEN_298; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_320 = io_in_14_valid ? io_in_14_bits_waddr : _GEN_301; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_324 = io_in_13_valid ? io_in_13_bits_len : _GEN_305; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_325 = io_in_13_valid ? io_in_13_bits_size : _GEN_306; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_327 = io_in_13_valid ? io_in_13_bits_mask : _GEN_308; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_328 = io_in_13_valid ? io_in_13_bits_data : _GEN_309; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_335 = io_in_13_valid ? io_in_13_bits_awid : _GEN_316; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_336 = io_in_13_valid ? io_in_13_bits_entryid : _GEN_317; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_339 = io_in_13_valid ? io_in_13_bits_waddr : _GEN_320; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_343 = io_in_12_valid ? io_in_12_bits_len : _GEN_324; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_344 = io_in_12_valid ? io_in_12_bits_size : _GEN_325; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_346 = io_in_12_valid ? io_in_12_bits_mask : _GEN_327; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_347 = io_in_12_valid ? io_in_12_bits_data : _GEN_328; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_354 = io_in_12_valid ? io_in_12_bits_awid : _GEN_335; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_355 = io_in_12_valid ? io_in_12_bits_entryid : _GEN_336; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_358 = io_in_12_valid ? io_in_12_bits_waddr : _GEN_339; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_362 = io_in_11_valid ? io_in_11_bits_len : _GEN_343; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_363 = io_in_11_valid ? io_in_11_bits_size : _GEN_344; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_365 = io_in_11_valid ? io_in_11_bits_mask : _GEN_346; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_366 = io_in_11_valid ? io_in_11_bits_data : _GEN_347; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_373 = io_in_11_valid ? io_in_11_bits_awid : _GEN_354; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_374 = io_in_11_valid ? io_in_11_bits_entryid : _GEN_355; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_377 = io_in_11_valid ? io_in_11_bits_waddr : _GEN_358; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_381 = io_in_10_valid ? io_in_10_bits_len : _GEN_362; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_382 = io_in_10_valid ? io_in_10_bits_size : _GEN_363; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_384 = io_in_10_valid ? io_in_10_bits_mask : _GEN_365; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_385 = io_in_10_valid ? io_in_10_bits_data : _GEN_366; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_392 = io_in_10_valid ? io_in_10_bits_awid : _GEN_373; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_393 = io_in_10_valid ? io_in_10_bits_entryid : _GEN_374; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_396 = io_in_10_valid ? io_in_10_bits_waddr : _GEN_377; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_400 = io_in_9_valid ? io_in_9_bits_len : _GEN_381; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_401 = io_in_9_valid ? io_in_9_bits_size : _GEN_382; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_403 = io_in_9_valid ? io_in_9_bits_mask : _GEN_384; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_404 = io_in_9_valid ? io_in_9_bits_data : _GEN_385; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_411 = io_in_9_valid ? io_in_9_bits_awid : _GEN_392; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_412 = io_in_9_valid ? io_in_9_bits_entryid : _GEN_393; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_415 = io_in_9_valid ? io_in_9_bits_waddr : _GEN_396; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_419 = io_in_8_valid ? io_in_8_bits_len : _GEN_400; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_420 = io_in_8_valid ? io_in_8_bits_size : _GEN_401; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_422 = io_in_8_valid ? io_in_8_bits_mask : _GEN_403; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_423 = io_in_8_valid ? io_in_8_bits_data : _GEN_404; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_430 = io_in_8_valid ? io_in_8_bits_awid : _GEN_411; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_431 = io_in_8_valid ? io_in_8_bits_entryid : _GEN_412; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_434 = io_in_8_valid ? io_in_8_bits_waddr : _GEN_415; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_438 = io_in_7_valid ? io_in_7_bits_len : _GEN_419; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_439 = io_in_7_valid ? io_in_7_bits_size : _GEN_420; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_441 = io_in_7_valid ? io_in_7_bits_mask : _GEN_422; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_442 = io_in_7_valid ? io_in_7_bits_data : _GEN_423; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_449 = io_in_7_valid ? io_in_7_bits_awid : _GEN_430; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_450 = io_in_7_valid ? io_in_7_bits_entryid : _GEN_431; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_453 = io_in_7_valid ? io_in_7_bits_waddr : _GEN_434; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_457 = io_in_6_valid ? io_in_6_bits_len : _GEN_438; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_458 = io_in_6_valid ? io_in_6_bits_size : _GEN_439; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_460 = io_in_6_valid ? io_in_6_bits_mask : _GEN_441; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_461 = io_in_6_valid ? io_in_6_bits_data : _GEN_442; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_468 = io_in_6_valid ? io_in_6_bits_awid : _GEN_449; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_469 = io_in_6_valid ? io_in_6_bits_entryid : _GEN_450; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_472 = io_in_6_valid ? io_in_6_bits_waddr : _GEN_453; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_476 = io_in_5_valid ? io_in_5_bits_len : _GEN_457; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_477 = io_in_5_valid ? io_in_5_bits_size : _GEN_458; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_479 = io_in_5_valid ? io_in_5_bits_mask : _GEN_460; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_480 = io_in_5_valid ? io_in_5_bits_data : _GEN_461; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_487 = io_in_5_valid ? io_in_5_bits_awid : _GEN_468; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_488 = io_in_5_valid ? io_in_5_bits_entryid : _GEN_469; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_491 = io_in_5_valid ? io_in_5_bits_waddr : _GEN_472; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_495 = io_in_4_valid ? io_in_4_bits_len : _GEN_476; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_496 = io_in_4_valid ? io_in_4_bits_size : _GEN_477; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_498 = io_in_4_valid ? io_in_4_bits_mask : _GEN_479; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_499 = io_in_4_valid ? io_in_4_bits_data : _GEN_480; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_506 = io_in_4_valid ? io_in_4_bits_awid : _GEN_487; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_507 = io_in_4_valid ? io_in_4_bits_entryid : _GEN_488; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_510 = io_in_4_valid ? io_in_4_bits_waddr : _GEN_491; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_514 = io_in_3_valid ? io_in_3_bits_len : _GEN_495; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_515 = io_in_3_valid ? io_in_3_bits_size : _GEN_496; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_517 = io_in_3_valid ? io_in_3_bits_mask : _GEN_498; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_518 = io_in_3_valid ? io_in_3_bits_data : _GEN_499; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_525 = io_in_3_valid ? io_in_3_bits_awid : _GEN_506; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_526 = io_in_3_valid ? io_in_3_bits_entryid : _GEN_507; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_529 = io_in_3_valid ? io_in_3_bits_waddr : _GEN_510; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_533 = io_in_2_valid ? io_in_2_bits_len : _GEN_514; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_534 = io_in_2_valid ? io_in_2_bits_size : _GEN_515; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_536 = io_in_2_valid ? io_in_2_bits_mask : _GEN_517; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_537 = io_in_2_valid ? io_in_2_bits_data : _GEN_518; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_544 = io_in_2_valid ? io_in_2_bits_awid : _GEN_525; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_545 = io_in_2_valid ? io_in_2_bits_entryid : _GEN_526; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_548 = io_in_2_valid ? io_in_2_bits_waddr : _GEN_529; // @[Arbiter.scala 141:26 143:19]
  wire [7:0] _GEN_552 = io_in_1_valid ? io_in_1_bits_len : _GEN_533; // @[Arbiter.scala 141:26 143:19]
  wire [2:0] _GEN_553 = io_in_1_valid ? io_in_1_bits_size : _GEN_534; // @[Arbiter.scala 141:26 143:19]
  wire [31:0] _GEN_555 = io_in_1_valid ? io_in_1_bits_mask : _GEN_536; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_556 = io_in_1_valid ? io_in_1_bits_data : _GEN_537; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_563 = io_in_1_valid ? io_in_1_bits_awid : _GEN_544; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_564 = io_in_1_valid ? io_in_1_bits_entryid : _GEN_545; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_567 = io_in_1_valid ? io_in_1_bits_waddr : _GEN_548; // @[Arbiter.scala 141:26 143:19]
  wire  _grant_T_29 = io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid | io_in_5_valid |
    io_in_6_valid | io_in_7_valid | io_in_8_valid | io_in_9_valid | io_in_10_valid | io_in_11_valid | io_in_12_valid |
    io_in_13_valid | io_in_14_valid | io_in_15_valid | io_in_16_valid | io_in_17_valid | io_in_18_valid | io_in_19_valid
     | io_in_20_valid | io_in_21_valid | io_in_22_valid | io_in_23_valid | io_in_24_valid | io_in_25_valid |
    io_in_26_valid | io_in_27_valid | io_in_28_valid | io_in_29_valid | io_in_30_valid; // @[Arbiter.scala 46:68]
  wire  grant_31 = ~_grant_T_29; // @[Arbiter.scala 46:78]
  assign io_out_valid = ~grant_31 | io_in_31_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_waddr = io_in_0_valid ? io_in_0_bits_waddr : _GEN_567; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_entryid = io_in_0_valid ? io_in_0_bits_entryid : _GEN_564; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_awid = io_in_0_valid ? io_in_0_bits_awid : _GEN_563; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_data = io_in_0_valid ? io_in_0_bits_data : _GEN_556; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_mask = io_in_0_valid ? io_in_0_bits_mask : _GEN_555; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : _GEN_553; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_len = io_in_0_valid ? io_in_0_bits_len : _GEN_552; // @[Arbiter.scala 141:26 143:19]
endmodule
module WriteStack(
  input          clock,
  input          reset,
  output         io_axiWriteReq_in_aw_ready,
  input          io_axiWriteReq_in_aw_valid,
  input  [13:0]  io_axiWriteReq_in_aw_bits_id,
  input  [34:0]  io_axiWriteReq_in_aw_bits_addr,
  input  [7:0]   io_axiWriteReq_in_aw_bits_len,
  input  [2:0]   io_axiWriteReq_in_aw_bits_size,
  input  [1:0]   io_axiWriteReq_in_aw_bits_burst,
  input          io_axiWriteReq_in_aw_bits_lock,
  input  [3:0]   io_axiWriteReq_in_aw_bits_cache,
  input  [2:0]   io_axiWriteReq_in_aw_bits_prot,
  input  [3:0]   io_axiWriteReq_in_aw_bits_qos,
  output         io_axiWriteReq_in_w_ready,
  input          io_axiWriteReq_in_w_valid,
  input  [255:0] io_axiWriteReq_in_w_bits_data,
  input  [31:0]  io_axiWriteReq_in_w_bits_strb,
  input          io_axiWriteReq_in_w_bits_last,
  input          io_axiMenWriteReq_out_aw_ready,
  output         io_axiMenWriteReq_out_aw_valid,
  output [13:0]  io_axiMenWriteReq_out_aw_bits_id,
  output [34:0]  io_axiMenWriteReq_out_aw_bits_addr,
  output [7:0]   io_axiMenWriteReq_out_aw_bits_len,
  output [2:0]   io_axiMenWriteReq_out_aw_bits_size,
  output [1:0]   io_axiMenWriteReq_out_aw_bits_burst,
  output         io_axiMenWriteReq_out_aw_bits_lock,
  output [3:0]   io_axiMenWriteReq_out_aw_bits_cache,
  output [2:0]   io_axiMenWriteReq_out_aw_bits_prot,
  output [3:0]   io_axiMenWriteReq_out_aw_bits_qos,
  input          io_axiMenWriteReq_out_w_ready,
  output         io_axiMenWriteReq_out_w_valid,
  output [255:0] io_axiMenWriteReq_out_w_bits_data,
  output [31:0]  io_axiMenWriteReq_out_w_bits_strb,
  output         io_axiMenWriteReq_out_w_bits_last,
  output         io_axiMenWriteResp_in_b_ready,
  input          io_axiMenWriteResp_in_b_valid,
  input  [13:0]  io_axiMenWriteResp_in_b_bits_id,
  input  [1:0]   io_axiMenWriteResp_in_b_bits_resp,
  input          io_axiWriteResp_out_b_ready,
  output         io_axiWriteResp_out_b_valid,
  output [13:0]  io_axiWriteResp_out_b_bits_id,
  output [1:0]   io_axiWriteResp_out_b_bits_resp,
  input          io_validReq_in_ready,
  output         io_validReq_in_valid,
  output [34:0]  io_validReq_in_bits_addr,
  output [18:0]  io_validReq_in_bits_source,
  output         io_validResp_out_ready,
  input          io_validResp_out_valid,
  input  [18:0]  io_validResp_out_bits_source,
  input          io_validResp_out_bits_validStatus
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [255:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [255:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [63:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [255:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [63:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [255:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [63:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [255:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [63:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [255:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [63:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [255:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [63:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [255:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [63:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [255:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [255:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [63:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [255:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [63:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [255:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [63:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [255:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [63:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [255:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [63:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [255:0] _RAND_203;
  reg [31:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [63:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [31:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [31:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [255:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [31:0] _RAND_221;
  reg [63:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [31:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [255:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [31:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [31:0] _RAND_234;
  reg [63:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [31:0] _RAND_241;
  reg [255:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [31:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [63:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [31:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [31:0] _RAND_254;
  reg [255:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [31:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [255:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [31:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [63:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [255:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [31:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [63:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [31:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [255:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [63:0] _RAND_300;
  reg [31:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [31:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [255:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [31:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [63:0] _RAND_313;
  reg [31:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
  reg [255:0] _RAND_320;
  reg [31:0] _RAND_321;
  reg [31:0] _RAND_322;
  reg [31:0] _RAND_323;
  reg [31:0] _RAND_324;
  reg [31:0] _RAND_325;
  reg [63:0] _RAND_326;
  reg [31:0] _RAND_327;
  reg [31:0] _RAND_328;
  reg [31:0] _RAND_329;
  reg [31:0] _RAND_330;
  reg [31:0] _RAND_331;
  reg [31:0] _RAND_332;
  reg [255:0] _RAND_333;
  reg [31:0] _RAND_334;
  reg [31:0] _RAND_335;
  reg [31:0] _RAND_336;
  reg [31:0] _RAND_337;
  reg [31:0] _RAND_338;
  reg [63:0] _RAND_339;
  reg [31:0] _RAND_340;
  reg [31:0] _RAND_341;
  reg [31:0] _RAND_342;
  reg [31:0] _RAND_343;
  reg [31:0] _RAND_344;
  reg [31:0] _RAND_345;
  reg [255:0] _RAND_346;
  reg [31:0] _RAND_347;
  reg [31:0] _RAND_348;
  reg [31:0] _RAND_349;
  reg [31:0] _RAND_350;
  reg [31:0] _RAND_351;
  reg [63:0] _RAND_352;
  reg [31:0] _RAND_353;
  reg [31:0] _RAND_354;
  reg [31:0] _RAND_355;
  reg [31:0] _RAND_356;
  reg [31:0] _RAND_357;
  reg [31:0] _RAND_358;
  reg [255:0] _RAND_359;
  reg [31:0] _RAND_360;
  reg [31:0] _RAND_361;
  reg [31:0] _RAND_362;
  reg [31:0] _RAND_363;
  reg [31:0] _RAND_364;
  reg [63:0] _RAND_365;
  reg [31:0] _RAND_366;
  reg [31:0] _RAND_367;
  reg [31:0] _RAND_368;
  reg [31:0] _RAND_369;
  reg [31:0] _RAND_370;
  reg [31:0] _RAND_371;
  reg [255:0] _RAND_372;
  reg [31:0] _RAND_373;
  reg [31:0] _RAND_374;
  reg [31:0] _RAND_375;
  reg [31:0] _RAND_376;
  reg [31:0] _RAND_377;
  reg [63:0] _RAND_378;
  reg [31:0] _RAND_379;
  reg [31:0] _RAND_380;
  reg [31:0] _RAND_381;
  reg [31:0] _RAND_382;
  reg [31:0] _RAND_383;
  reg [31:0] _RAND_384;
  reg [255:0] _RAND_385;
  reg [31:0] _RAND_386;
  reg [31:0] _RAND_387;
  reg [31:0] _RAND_388;
  reg [31:0] _RAND_389;
  reg [31:0] _RAND_390;
  reg [63:0] _RAND_391;
  reg [31:0] _RAND_392;
  reg [31:0] _RAND_393;
  reg [31:0] _RAND_394;
  reg [31:0] _RAND_395;
  reg [31:0] _RAND_396;
  reg [31:0] _RAND_397;
  reg [255:0] _RAND_398;
  reg [31:0] _RAND_399;
  reg [31:0] _RAND_400;
  reg [31:0] _RAND_401;
  reg [31:0] _RAND_402;
  reg [31:0] _RAND_403;
  reg [63:0] _RAND_404;
  reg [31:0] _RAND_405;
  reg [31:0] _RAND_406;
  reg [31:0] _RAND_407;
  reg [31:0] _RAND_408;
  reg [31:0] _RAND_409;
  reg [31:0] _RAND_410;
  reg [255:0] _RAND_411;
  reg [31:0] _RAND_412;
  reg [31:0] _RAND_413;
  reg [31:0] _RAND_414;
  reg [31:0] _RAND_415;
`endif // RANDOMIZE_REG_INIT
  wire  wreqArb_io_in_0_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_0_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_0_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_0_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_0_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_0_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_0_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_0_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_1_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_1_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_1_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_1_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_1_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_1_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_1_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_1_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_2_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_2_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_2_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_2_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_2_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_2_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_2_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_2_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_3_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_3_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_3_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_3_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_3_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_3_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_3_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_3_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_4_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_4_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_4_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_4_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_4_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_4_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_4_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_4_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_5_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_5_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_5_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_5_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_5_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_5_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_5_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_5_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_6_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_6_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_6_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_6_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_6_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_6_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_6_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_6_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_7_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_7_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_7_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_7_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_7_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_7_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_7_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_7_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_8_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_8_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_8_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_8_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_8_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_8_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_8_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_8_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_9_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_9_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_9_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_9_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_9_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_9_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_9_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_9_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_10_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_10_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_10_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_10_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_10_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_10_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_10_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_10_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_11_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_11_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_11_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_11_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_11_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_11_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_11_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_11_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_12_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_12_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_12_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_12_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_12_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_12_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_12_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_12_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_13_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_13_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_13_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_13_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_13_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_13_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_13_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_13_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_14_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_14_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_14_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_14_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_14_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_14_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_14_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_14_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_15_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_15_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_15_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_15_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_15_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_15_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_15_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_15_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_16_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_16_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_16_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_16_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_16_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_16_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_16_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_16_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_17_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_17_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_17_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_17_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_17_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_17_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_17_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_17_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_18_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_18_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_18_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_18_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_18_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_18_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_18_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_18_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_19_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_19_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_19_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_19_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_19_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_19_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_19_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_19_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_20_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_20_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_20_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_20_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_20_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_20_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_20_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_20_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_21_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_21_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_21_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_21_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_21_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_21_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_21_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_21_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_22_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_22_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_22_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_22_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_22_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_22_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_22_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_22_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_23_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_23_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_23_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_23_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_23_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_23_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_23_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_23_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_24_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_24_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_24_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_24_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_24_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_24_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_24_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_24_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_25_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_25_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_25_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_25_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_25_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_25_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_25_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_25_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_26_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_26_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_26_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_26_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_26_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_26_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_26_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_26_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_27_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_27_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_27_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_27_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_27_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_27_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_27_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_27_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_28_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_28_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_28_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_28_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_28_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_28_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_28_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_28_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_29_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_29_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_29_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_29_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_29_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_29_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_29_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_29_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_30_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_30_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_30_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_30_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_30_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_30_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_30_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_30_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_in_31_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_in_31_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_in_31_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_in_31_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_in_31_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_in_31_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_in_31_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_in_31_bits_len; // @[WriteStack.scala 60:23]
  wire  wreqArb_io_out_valid; // @[WriteStack.scala 60:23]
  wire [34:0] wreqArb_io_out_bits_waddr; // @[WriteStack.scala 60:23]
  wire [4:0] wreqArb_io_out_bits_entryid; // @[WriteStack.scala 60:23]
  wire [13:0] wreqArb_io_out_bits_awid; // @[WriteStack.scala 60:23]
  wire [255:0] wreqArb_io_out_bits_data; // @[WriteStack.scala 60:23]
  wire [31:0] wreqArb_io_out_bits_mask; // @[WriteStack.scala 60:23]
  wire [2:0] wreqArb_io_out_bits_size; // @[WriteStack.scala 60:23]
  wire [7:0] wreqArb_io_out_bits_len; // @[WriteStack.scala 60:23]
  wire  awreqArb_io_in_0_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_0_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_0_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_0_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_0_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_0_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_0_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_0_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_1_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_1_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_1_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_1_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_1_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_1_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_1_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_1_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_2_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_2_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_2_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_2_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_2_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_2_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_2_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_2_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_3_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_3_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_3_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_3_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_3_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_3_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_3_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_3_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_4_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_4_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_4_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_4_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_4_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_4_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_4_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_4_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_5_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_5_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_5_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_5_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_5_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_5_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_5_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_5_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_6_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_6_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_6_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_6_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_6_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_6_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_6_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_6_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_7_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_7_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_7_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_7_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_7_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_7_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_7_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_7_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_8_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_8_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_8_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_8_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_8_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_8_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_8_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_8_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_9_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_9_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_9_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_9_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_9_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_9_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_9_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_9_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_10_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_10_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_10_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_10_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_10_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_10_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_10_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_10_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_11_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_11_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_11_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_11_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_11_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_11_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_11_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_11_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_12_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_12_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_12_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_12_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_12_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_12_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_12_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_12_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_13_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_13_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_13_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_13_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_13_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_13_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_13_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_13_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_14_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_14_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_14_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_14_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_14_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_14_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_14_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_14_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_15_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_15_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_15_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_15_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_15_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_15_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_15_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_15_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_16_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_16_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_16_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_16_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_16_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_16_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_16_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_16_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_17_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_17_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_17_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_17_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_17_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_17_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_17_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_17_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_18_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_18_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_18_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_18_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_18_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_18_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_18_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_18_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_19_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_19_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_19_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_19_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_19_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_19_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_19_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_19_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_20_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_20_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_20_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_20_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_20_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_20_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_20_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_20_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_21_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_21_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_21_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_21_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_21_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_21_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_21_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_21_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_22_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_22_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_22_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_22_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_22_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_22_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_22_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_22_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_23_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_23_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_23_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_23_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_23_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_23_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_23_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_23_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_24_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_24_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_24_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_24_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_24_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_24_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_24_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_24_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_25_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_25_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_25_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_25_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_25_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_25_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_25_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_25_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_26_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_26_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_26_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_26_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_26_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_26_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_26_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_26_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_27_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_27_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_27_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_27_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_27_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_27_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_27_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_27_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_28_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_28_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_28_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_28_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_28_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_28_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_28_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_28_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_29_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_29_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_29_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_29_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_29_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_29_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_29_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_29_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_30_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_30_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_30_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_30_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_30_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_30_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_30_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_30_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_in_31_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_in_31_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_in_31_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_in_31_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_in_31_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_in_31_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_in_31_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_in_31_bits_len; // @[WriteStack.scala 61:24]
  wire  awreqArb_io_out_valid; // @[WriteStack.scala 61:24]
  wire [34:0] awreqArb_io_out_bits_waddr; // @[WriteStack.scala 61:24]
  wire [4:0] awreqArb_io_out_bits_entryid; // @[WriteStack.scala 61:24]
  wire [13:0] awreqArb_io_out_bits_awid; // @[WriteStack.scala 61:24]
  wire [255:0] awreqArb_io_out_bits_data; // @[WriteStack.scala 61:24]
  wire [31:0] awreqArb_io_out_bits_mask; // @[WriteStack.scala 61:24]
  wire [2:0] awreqArb_io_out_bits_size; // @[WriteStack.scala 61:24]
  wire [7:0] awreqArb_io_out_bits_len; // @[WriteStack.scala 61:24]
  wire  validreqArb_io_in_0_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_0_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_0_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_0_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_0_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_0_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_0_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_0_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_1_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_1_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_1_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_1_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_1_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_1_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_1_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_1_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_2_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_2_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_2_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_2_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_2_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_2_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_2_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_2_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_3_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_3_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_3_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_3_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_3_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_3_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_3_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_3_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_4_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_4_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_4_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_4_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_4_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_4_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_4_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_4_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_5_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_5_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_5_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_5_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_5_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_5_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_5_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_5_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_6_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_6_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_6_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_6_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_6_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_6_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_6_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_6_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_7_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_7_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_7_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_7_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_7_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_7_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_7_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_7_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_8_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_8_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_8_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_8_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_8_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_8_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_8_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_8_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_9_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_9_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_9_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_9_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_9_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_9_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_9_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_9_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_10_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_10_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_10_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_10_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_10_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_10_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_10_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_10_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_11_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_11_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_11_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_11_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_11_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_11_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_11_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_11_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_12_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_12_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_12_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_12_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_12_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_12_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_12_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_12_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_13_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_13_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_13_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_13_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_13_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_13_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_13_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_13_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_14_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_14_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_14_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_14_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_14_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_14_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_14_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_14_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_15_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_15_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_15_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_15_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_15_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_15_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_15_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_15_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_16_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_16_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_16_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_16_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_16_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_16_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_16_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_16_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_17_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_17_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_17_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_17_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_17_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_17_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_17_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_17_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_18_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_18_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_18_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_18_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_18_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_18_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_18_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_18_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_19_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_19_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_19_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_19_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_19_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_19_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_19_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_19_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_20_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_20_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_20_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_20_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_20_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_20_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_20_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_20_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_21_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_21_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_21_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_21_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_21_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_21_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_21_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_21_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_22_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_22_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_22_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_22_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_22_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_22_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_22_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_22_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_23_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_23_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_23_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_23_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_23_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_23_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_23_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_23_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_24_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_24_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_24_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_24_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_24_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_24_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_24_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_24_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_25_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_25_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_25_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_25_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_25_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_25_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_25_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_25_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_26_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_26_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_26_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_26_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_26_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_26_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_26_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_26_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_27_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_27_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_27_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_27_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_27_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_27_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_27_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_27_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_28_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_28_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_28_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_28_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_28_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_28_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_28_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_28_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_29_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_29_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_29_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_29_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_29_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_29_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_29_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_29_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_30_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_30_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_30_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_30_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_30_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_30_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_30_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_30_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_in_31_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_in_31_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_in_31_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_in_31_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_in_31_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_in_31_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_in_31_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_in_31_bits_len; // @[WriteStack.scala 62:27]
  wire  validreqArb_io_out_valid; // @[WriteStack.scala 62:27]
  wire [34:0] validreqArb_io_out_bits_waddr; // @[WriteStack.scala 62:27]
  wire [4:0] validreqArb_io_out_bits_entryid; // @[WriteStack.scala 62:27]
  wire [13:0] validreqArb_io_out_bits_awid; // @[WriteStack.scala 62:27]
  wire [255:0] validreqArb_io_out_bits_data; // @[WriteStack.scala 62:27]
  wire [31:0] validreqArb_io_out_bits_mask; // @[WriteStack.scala 62:27]
  wire [2:0] validreqArb_io_out_bits_size; // @[WriteStack.scala 62:27]
  wire [7:0] validreqArb_io_out_bits_len; // @[WriteStack.scala 62:27]
  reg  writeStack_0_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_0_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_0_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_0_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_0_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_0_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_0_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_0_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_0_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_0_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_0_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_0_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_0_len; // @[WriteStack.scala 56:27]
  reg  writeStack_1_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_1_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_1_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_1_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_1_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_1_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_1_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_1_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_1_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_1_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_1_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_1_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_1_len; // @[WriteStack.scala 56:27]
  reg  writeStack_2_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_2_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_2_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_2_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_2_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_2_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_2_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_2_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_2_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_2_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_2_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_2_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_2_len; // @[WriteStack.scala 56:27]
  reg  writeStack_3_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_3_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_3_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_3_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_3_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_3_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_3_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_3_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_3_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_3_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_3_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_3_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_3_len; // @[WriteStack.scala 56:27]
  reg  writeStack_4_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_4_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_4_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_4_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_4_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_4_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_4_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_4_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_4_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_4_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_4_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_4_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_4_len; // @[WriteStack.scala 56:27]
  reg  writeStack_5_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_5_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_5_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_5_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_5_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_5_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_5_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_5_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_5_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_5_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_5_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_5_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_5_len; // @[WriteStack.scala 56:27]
  reg  writeStack_6_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_6_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_6_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_6_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_6_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_6_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_6_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_6_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_6_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_6_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_6_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_6_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_6_len; // @[WriteStack.scala 56:27]
  reg  writeStack_7_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_7_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_7_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_7_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_7_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_7_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_7_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_7_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_7_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_7_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_7_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_7_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_7_len; // @[WriteStack.scala 56:27]
  reg  writeStack_8_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_8_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_8_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_8_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_8_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_8_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_8_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_8_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_8_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_8_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_8_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_8_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_8_len; // @[WriteStack.scala 56:27]
  reg  writeStack_9_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_9_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_9_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_9_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_9_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_9_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_9_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_9_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_9_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_9_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_9_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_9_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_9_len; // @[WriteStack.scala 56:27]
  reg  writeStack_10_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_10_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_10_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_10_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_10_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_10_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_10_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_10_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_10_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_10_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_10_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_10_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_10_len; // @[WriteStack.scala 56:27]
  reg  writeStack_11_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_11_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_11_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_11_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_11_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_11_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_11_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_11_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_11_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_11_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_11_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_11_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_11_len; // @[WriteStack.scala 56:27]
  reg  writeStack_12_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_12_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_12_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_12_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_12_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_12_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_12_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_12_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_12_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_12_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_12_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_12_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_12_len; // @[WriteStack.scala 56:27]
  reg  writeStack_13_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_13_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_13_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_13_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_13_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_13_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_13_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_13_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_13_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_13_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_13_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_13_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_13_len; // @[WriteStack.scala 56:27]
  reg  writeStack_14_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_14_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_14_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_14_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_14_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_14_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_14_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_14_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_14_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_14_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_14_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_14_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_14_len; // @[WriteStack.scala 56:27]
  reg  writeStack_15_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_15_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_15_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_15_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_15_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_15_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_15_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_15_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_15_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_15_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_15_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_15_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_15_len; // @[WriteStack.scala 56:27]
  reg  writeStack_16_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_16_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_16_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_16_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_16_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_16_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_16_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_16_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_16_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_16_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_16_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_16_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_16_len; // @[WriteStack.scala 56:27]
  reg  writeStack_17_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_17_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_17_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_17_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_17_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_17_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_17_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_17_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_17_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_17_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_17_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_17_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_17_len; // @[WriteStack.scala 56:27]
  reg  writeStack_18_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_18_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_18_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_18_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_18_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_18_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_18_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_18_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_18_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_18_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_18_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_18_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_18_len; // @[WriteStack.scala 56:27]
  reg  writeStack_19_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_19_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_19_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_19_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_19_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_19_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_19_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_19_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_19_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_19_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_19_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_19_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_19_len; // @[WriteStack.scala 56:27]
  reg  writeStack_20_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_20_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_20_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_20_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_20_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_20_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_20_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_20_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_20_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_20_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_20_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_20_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_20_len; // @[WriteStack.scala 56:27]
  reg  writeStack_21_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_21_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_21_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_21_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_21_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_21_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_21_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_21_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_21_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_21_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_21_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_21_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_21_len; // @[WriteStack.scala 56:27]
  reg  writeStack_22_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_22_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_22_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_22_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_22_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_22_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_22_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_22_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_22_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_22_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_22_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_22_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_22_len; // @[WriteStack.scala 56:27]
  reg  writeStack_23_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_23_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_23_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_23_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_23_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_23_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_23_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_23_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_23_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_23_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_23_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_23_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_23_len; // @[WriteStack.scala 56:27]
  reg  writeStack_24_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_24_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_24_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_24_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_24_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_24_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_24_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_24_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_24_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_24_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_24_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_24_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_24_len; // @[WriteStack.scala 56:27]
  reg  writeStack_25_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_25_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_25_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_25_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_25_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_25_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_25_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_25_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_25_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_25_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_25_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_25_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_25_len; // @[WriteStack.scala 56:27]
  reg  writeStack_26_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_26_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_26_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_26_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_26_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_26_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_26_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_26_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_26_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_26_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_26_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_26_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_26_len; // @[WriteStack.scala 56:27]
  reg  writeStack_27_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_27_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_27_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_27_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_27_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_27_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_27_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_27_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_27_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_27_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_27_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_27_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_27_len; // @[WriteStack.scala 56:27]
  reg  writeStack_28_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_28_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_28_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_28_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_28_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_28_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_28_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_28_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_28_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_28_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_28_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_28_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_28_len; // @[WriteStack.scala 56:27]
  reg  writeStack_29_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_29_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_29_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_29_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_29_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_29_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_29_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_29_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_29_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_29_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_29_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_29_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_29_len; // @[WriteStack.scala 56:27]
  reg  writeStack_30_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_30_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_30_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_30_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_30_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_30_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_30_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_30_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_30_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_30_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_30_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_30_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_30_len; // @[WriteStack.scala 56:27]
  reg  writeStack_31_wvalid; // @[WriteStack.scala 56:27]
  reg [34:0] writeStack_31_waddr; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_31_wstatus; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_31_entryid; // @[WriteStack.scala 56:27]
  reg [13:0] writeStack_31_awid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_31_entryFifoid; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_31_validFifoId; // @[WriteStack.scala 56:27]
  reg [4:0] writeStack_31_waitWFifoId; // @[WriteStack.scala 56:27]
  reg [255:0] writeStack_31_data; // @[WriteStack.scala 56:27]
  reg [31:0] writeStack_31_mask; // @[WriteStack.scala 56:27]
  reg [1:0] writeStack_31_validStatus; // @[WriteStack.scala 56:27]
  reg [2:0] writeStack_31_size; // @[WriteStack.scala 56:27]
  reg [7:0] writeStack_31_len; // @[WriteStack.scala 56:27]
  wire [7:0] full_lo_lo = {writeStack_24_wvalid,writeStack_25_wvalid,writeStack_26_wvalid,writeStack_27_wvalid,
    writeStack_28_wvalid,writeStack_29_wvalid,writeStack_30_wvalid,writeStack_31_wvalid}; // @[Cat.scala 31:58]
  wire [15:0] full_lo = {writeStack_16_wvalid,writeStack_17_wvalid,writeStack_18_wvalid,writeStack_19_wvalid,
    writeStack_20_wvalid,writeStack_21_wvalid,writeStack_22_wvalid,writeStack_23_wvalid,full_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] full_hi_lo = {writeStack_8_wvalid,writeStack_9_wvalid,writeStack_10_wvalid,writeStack_11_wvalid,
    writeStack_12_wvalid,writeStack_13_wvalid,writeStack_14_wvalid,writeStack_15_wvalid}; // @[Cat.scala 31:58]
  wire [31:0] _full_T = {writeStack_0_wvalid,writeStack_1_wvalid,writeStack_2_wvalid,writeStack_3_wvalid,
    writeStack_4_wvalid,writeStack_5_wvalid,writeStack_6_wvalid,writeStack_7_wvalid,full_hi_lo,full_lo}; // @[Cat.scala 31:58]
  wire  full = &_full_T; // @[WriteStack.scala 65:44]
  wire  alloc = ~full & io_axiWriteReq_in_aw_valid; // @[WriteStack.scala 66:21]
  wire  _idxInsert_T = ~writeStack_0_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_1 = ~writeStack_1_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_2 = ~writeStack_2_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_3 = ~writeStack_3_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_4 = ~writeStack_4_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_5 = ~writeStack_5_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_6 = ~writeStack_6_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_7 = ~writeStack_7_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_8 = ~writeStack_8_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_9 = ~writeStack_9_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_10 = ~writeStack_10_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_11 = ~writeStack_11_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_12 = ~writeStack_12_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_13 = ~writeStack_13_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_14 = ~writeStack_14_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_15 = ~writeStack_15_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_16 = ~writeStack_16_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_17 = ~writeStack_17_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_18 = ~writeStack_18_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_19 = ~writeStack_19_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_20 = ~writeStack_20_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_21 = ~writeStack_21_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_22 = ~writeStack_22_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_23 = ~writeStack_23_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_24 = ~writeStack_24_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_25 = ~writeStack_25_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_26 = ~writeStack_26_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_27 = ~writeStack_27_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_28 = ~writeStack_28_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_29 = ~writeStack_29_wvalid; // @[WriteStack.scala 68:60]
  wire  _idxInsert_T_30 = ~writeStack_30_wvalid; // @[WriteStack.scala 68:60]
  wire [4:0] _idxInsert_T_32 = _idxInsert_T_30 ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_33 = _idxInsert_T_29 ? 5'h1d : _idxInsert_T_32; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_34 = _idxInsert_T_28 ? 5'h1c : _idxInsert_T_33; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_35 = _idxInsert_T_27 ? 5'h1b : _idxInsert_T_34; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_36 = _idxInsert_T_26 ? 5'h1a : _idxInsert_T_35; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_37 = _idxInsert_T_25 ? 5'h19 : _idxInsert_T_36; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_38 = _idxInsert_T_24 ? 5'h18 : _idxInsert_T_37; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_39 = _idxInsert_T_23 ? 5'h17 : _idxInsert_T_38; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_40 = _idxInsert_T_22 ? 5'h16 : _idxInsert_T_39; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_41 = _idxInsert_T_21 ? 5'h15 : _idxInsert_T_40; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_42 = _idxInsert_T_20 ? 5'h14 : _idxInsert_T_41; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_43 = _idxInsert_T_19 ? 5'h13 : _idxInsert_T_42; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_44 = _idxInsert_T_18 ? 5'h12 : _idxInsert_T_43; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_45 = _idxInsert_T_17 ? 5'h11 : _idxInsert_T_44; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_46 = _idxInsert_T_16 ? 5'h10 : _idxInsert_T_45; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_47 = _idxInsert_T_15 ? 5'hf : _idxInsert_T_46; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_48 = _idxInsert_T_14 ? 5'he : _idxInsert_T_47; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_49 = _idxInsert_T_13 ? 5'hd : _idxInsert_T_48; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_50 = _idxInsert_T_12 ? 5'hc : _idxInsert_T_49; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_51 = _idxInsert_T_11 ? 5'hb : _idxInsert_T_50; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_52 = _idxInsert_T_10 ? 5'ha : _idxInsert_T_51; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_53 = _idxInsert_T_9 ? 5'h9 : _idxInsert_T_52; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_54 = _idxInsert_T_8 ? 5'h8 : _idxInsert_T_53; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_55 = _idxInsert_T_7 ? 5'h7 : _idxInsert_T_54; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_56 = _idxInsert_T_6 ? 5'h6 : _idxInsert_T_55; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_57 = _idxInsert_T_5 ? 5'h5 : _idxInsert_T_56; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_58 = _idxInsert_T_4 ? 5'h4 : _idxInsert_T_57; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_59 = _idxInsert_T_3 ? 5'h3 : _idxInsert_T_58; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_60 = _idxInsert_T_2 ? 5'h2 : _idxInsert_T_59; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_61 = _idxInsert_T_1 ? 5'h1 : _idxInsert_T_60; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_62 = _idxInsert_T ? 5'h0 : _idxInsert_T_61; // @[Mux.scala 47:70]
  wire [4:0] idxInsert = alloc ? _idxInsert_T_62 : 5'h0; // @[WriteStack.scala 68:22]
  wire  _GEN_0 = 5'h0 == idxInsert | writeStack_0_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_1 = 5'h1 == idxInsert | writeStack_1_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_2 = 5'h2 == idxInsert | writeStack_2_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_3 = 5'h3 == idxInsert | writeStack_3_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_4 = 5'h4 == idxInsert | writeStack_4_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_5 = 5'h5 == idxInsert | writeStack_5_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_6 = 5'h6 == idxInsert | writeStack_6_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_7 = 5'h7 == idxInsert | writeStack_7_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_8 = 5'h8 == idxInsert | writeStack_8_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_9 = 5'h9 == idxInsert | writeStack_9_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_10 = 5'ha == idxInsert | writeStack_10_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_11 = 5'hb == idxInsert | writeStack_11_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_12 = 5'hc == idxInsert | writeStack_12_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_13 = 5'hd == idxInsert | writeStack_13_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_14 = 5'he == idxInsert | writeStack_14_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_15 = 5'hf == idxInsert | writeStack_15_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_16 = 5'h10 == idxInsert | writeStack_16_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_17 = 5'h11 == idxInsert | writeStack_17_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_18 = 5'h12 == idxInsert | writeStack_18_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_19 = 5'h13 == idxInsert | writeStack_19_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_20 = 5'h14 == idxInsert | writeStack_20_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_21 = 5'h15 == idxInsert | writeStack_21_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_22 = 5'h16 == idxInsert | writeStack_22_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_23 = 5'h17 == idxInsert | writeStack_23_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_24 = 5'h18 == idxInsert | writeStack_24_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_25 = 5'h19 == idxInsert | writeStack_25_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_26 = 5'h1a == idxInsert | writeStack_26_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_27 = 5'h1b == idxInsert | writeStack_27_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_28 = 5'h1c == idxInsert | writeStack_28_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_29 = 5'h1d == idxInsert | writeStack_29_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_30 = 5'h1e == idxInsert | writeStack_30_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire  _GEN_31 = 5'h1f == idxInsert | writeStack_31_wvalid; // @[WriteStack.scala 73:{19,19} 56:27]
  wire [1:0] _GEN_64 = 5'h0 == idxInsert ? 2'h1 : writeStack_0_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_65 = 5'h1 == idxInsert ? 2'h1 : writeStack_1_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_66 = 5'h2 == idxInsert ? 2'h1 : writeStack_2_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_67 = 5'h3 == idxInsert ? 2'h1 : writeStack_3_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_68 = 5'h4 == idxInsert ? 2'h1 : writeStack_4_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_69 = 5'h5 == idxInsert ? 2'h1 : writeStack_5_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_70 = 5'h6 == idxInsert ? 2'h1 : writeStack_6_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_71 = 5'h7 == idxInsert ? 2'h1 : writeStack_7_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_72 = 5'h8 == idxInsert ? 2'h1 : writeStack_8_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_73 = 5'h9 == idxInsert ? 2'h1 : writeStack_9_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_74 = 5'ha == idxInsert ? 2'h1 : writeStack_10_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_75 = 5'hb == idxInsert ? 2'h1 : writeStack_11_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_76 = 5'hc == idxInsert ? 2'h1 : writeStack_12_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_77 = 5'hd == idxInsert ? 2'h1 : writeStack_13_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_78 = 5'he == idxInsert ? 2'h1 : writeStack_14_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_79 = 5'hf == idxInsert ? 2'h1 : writeStack_15_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_80 = 5'h10 == idxInsert ? 2'h1 : writeStack_16_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_81 = 5'h11 == idxInsert ? 2'h1 : writeStack_17_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_82 = 5'h12 == idxInsert ? 2'h1 : writeStack_18_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_83 = 5'h13 == idxInsert ? 2'h1 : writeStack_19_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_84 = 5'h14 == idxInsert ? 2'h1 : writeStack_20_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_85 = 5'h15 == idxInsert ? 2'h1 : writeStack_21_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_86 = 5'h16 == idxInsert ? 2'h1 : writeStack_22_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_87 = 5'h17 == idxInsert ? 2'h1 : writeStack_23_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_88 = 5'h18 == idxInsert ? 2'h1 : writeStack_24_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_89 = 5'h19 == idxInsert ? 2'h1 : writeStack_25_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_90 = 5'h1a == idxInsert ? 2'h1 : writeStack_26_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_91 = 5'h1b == idxInsert ? 2'h1 : writeStack_27_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_92 = 5'h1c == idxInsert ? 2'h1 : writeStack_28_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_93 = 5'h1d == idxInsert ? 2'h1 : writeStack_29_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_94 = 5'h1e == idxInsert ? 2'h1 : writeStack_30_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_95 = 5'h1f == idxInsert ? 2'h1 : writeStack_31_wstatus; // @[WriteStack.scala 75:{19,19} 56:27]
  wire [1:0] _GEN_96 = 5'h0 == idxInsert ? 2'h1 : writeStack_0_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_97 = 5'h1 == idxInsert ? 2'h1 : writeStack_1_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_98 = 5'h2 == idxInsert ? 2'h1 : writeStack_2_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_99 = 5'h3 == idxInsert ? 2'h1 : writeStack_3_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_100 = 5'h4 == idxInsert ? 2'h1 : writeStack_4_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_101 = 5'h5 == idxInsert ? 2'h1 : writeStack_5_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_102 = 5'h6 == idxInsert ? 2'h1 : writeStack_6_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_103 = 5'h7 == idxInsert ? 2'h1 : writeStack_7_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_104 = 5'h8 == idxInsert ? 2'h1 : writeStack_8_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_105 = 5'h9 == idxInsert ? 2'h1 : writeStack_9_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_106 = 5'ha == idxInsert ? 2'h1 : writeStack_10_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_107 = 5'hb == idxInsert ? 2'h1 : writeStack_11_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_108 = 5'hc == idxInsert ? 2'h1 : writeStack_12_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_109 = 5'hd == idxInsert ? 2'h1 : writeStack_13_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_110 = 5'he == idxInsert ? 2'h1 : writeStack_14_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_111 = 5'hf == idxInsert ? 2'h1 : writeStack_15_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_112 = 5'h10 == idxInsert ? 2'h1 : writeStack_16_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_113 = 5'h11 == idxInsert ? 2'h1 : writeStack_17_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_114 = 5'h12 == idxInsert ? 2'h1 : writeStack_18_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_115 = 5'h13 == idxInsert ? 2'h1 : writeStack_19_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_116 = 5'h14 == idxInsert ? 2'h1 : writeStack_20_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_117 = 5'h15 == idxInsert ? 2'h1 : writeStack_21_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_118 = 5'h16 == idxInsert ? 2'h1 : writeStack_22_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_119 = 5'h17 == idxInsert ? 2'h1 : writeStack_23_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_120 = 5'h18 == idxInsert ? 2'h1 : writeStack_24_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_121 = 5'h19 == idxInsert ? 2'h1 : writeStack_25_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_122 = 5'h1a == idxInsert ? 2'h1 : writeStack_26_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_123 = 5'h1b == idxInsert ? 2'h1 : writeStack_27_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_124 = 5'h1c == idxInsert ? 2'h1 : writeStack_28_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_125 = 5'h1d == idxInsert ? 2'h1 : writeStack_29_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_126 = 5'h1e == idxInsert ? 2'h1 : writeStack_30_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire [1:0] _GEN_127 = 5'h1f == idxInsert ? 2'h1 : writeStack_31_validStatus; // @[WriteStack.scala 76:{23,23} 56:27]
  wire  _GEN_288 = alloc ? _GEN_0 : writeStack_0_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_289 = alloc ? _GEN_1 : writeStack_1_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_290 = alloc ? _GEN_2 : writeStack_2_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_291 = alloc ? _GEN_3 : writeStack_3_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_292 = alloc ? _GEN_4 : writeStack_4_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_293 = alloc ? _GEN_5 : writeStack_5_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_294 = alloc ? _GEN_6 : writeStack_6_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_295 = alloc ? _GEN_7 : writeStack_7_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_296 = alloc ? _GEN_8 : writeStack_8_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_297 = alloc ? _GEN_9 : writeStack_9_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_298 = alloc ? _GEN_10 : writeStack_10_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_299 = alloc ? _GEN_11 : writeStack_11_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_300 = alloc ? _GEN_12 : writeStack_12_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_301 = alloc ? _GEN_13 : writeStack_13_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_302 = alloc ? _GEN_14 : writeStack_14_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_303 = alloc ? _GEN_15 : writeStack_15_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_304 = alloc ? _GEN_16 : writeStack_16_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_305 = alloc ? _GEN_17 : writeStack_17_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_306 = alloc ? _GEN_18 : writeStack_18_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_307 = alloc ? _GEN_19 : writeStack_19_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_308 = alloc ? _GEN_20 : writeStack_20_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_309 = alloc ? _GEN_21 : writeStack_21_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_310 = alloc ? _GEN_22 : writeStack_22_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_311 = alloc ? _GEN_23 : writeStack_23_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_312 = alloc ? _GEN_24 : writeStack_24_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_313 = alloc ? _GEN_25 : writeStack_25_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_314 = alloc ? _GEN_26 : writeStack_26_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_315 = alloc ? _GEN_27 : writeStack_27_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_316 = alloc ? _GEN_28 : writeStack_28_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_317 = alloc ? _GEN_29 : writeStack_29_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_318 = alloc ? _GEN_30 : writeStack_30_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire  _GEN_319 = alloc ? _GEN_31 : writeStack_31_wvalid; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_352 = alloc ? _GEN_64 : writeStack_0_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_353 = alloc ? _GEN_65 : writeStack_1_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_354 = alloc ? _GEN_66 : writeStack_2_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_355 = alloc ? _GEN_67 : writeStack_3_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_356 = alloc ? _GEN_68 : writeStack_4_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_357 = alloc ? _GEN_69 : writeStack_5_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_358 = alloc ? _GEN_70 : writeStack_6_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_359 = alloc ? _GEN_71 : writeStack_7_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_360 = alloc ? _GEN_72 : writeStack_8_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_361 = alloc ? _GEN_73 : writeStack_9_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_362 = alloc ? _GEN_74 : writeStack_10_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_363 = alloc ? _GEN_75 : writeStack_11_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_364 = alloc ? _GEN_76 : writeStack_12_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_365 = alloc ? _GEN_77 : writeStack_13_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_366 = alloc ? _GEN_78 : writeStack_14_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_367 = alloc ? _GEN_79 : writeStack_15_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_368 = alloc ? _GEN_80 : writeStack_16_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_369 = alloc ? _GEN_81 : writeStack_17_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_370 = alloc ? _GEN_82 : writeStack_18_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_371 = alloc ? _GEN_83 : writeStack_19_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_372 = alloc ? _GEN_84 : writeStack_20_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_373 = alloc ? _GEN_85 : writeStack_21_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_374 = alloc ? _GEN_86 : writeStack_22_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_375 = alloc ? _GEN_87 : writeStack_23_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_376 = alloc ? _GEN_88 : writeStack_24_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_377 = alloc ? _GEN_89 : writeStack_25_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_378 = alloc ? _GEN_90 : writeStack_26_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_379 = alloc ? _GEN_91 : writeStack_27_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_380 = alloc ? _GEN_92 : writeStack_28_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_381 = alloc ? _GEN_93 : writeStack_29_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_382 = alloc ? _GEN_94 : writeStack_30_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_383 = alloc ? _GEN_95 : writeStack_31_wstatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_384 = alloc ? _GEN_96 : writeStack_0_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_385 = alloc ? _GEN_97 : writeStack_1_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_386 = alloc ? _GEN_98 : writeStack_2_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_387 = alloc ? _GEN_99 : writeStack_3_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_388 = alloc ? _GEN_100 : writeStack_4_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_389 = alloc ? _GEN_101 : writeStack_5_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_390 = alloc ? _GEN_102 : writeStack_6_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_391 = alloc ? _GEN_103 : writeStack_7_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_392 = alloc ? _GEN_104 : writeStack_8_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_393 = alloc ? _GEN_105 : writeStack_9_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_394 = alloc ? _GEN_106 : writeStack_10_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_395 = alloc ? _GEN_107 : writeStack_11_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_396 = alloc ? _GEN_108 : writeStack_12_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_397 = alloc ? _GEN_109 : writeStack_13_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_398 = alloc ? _GEN_110 : writeStack_14_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_399 = alloc ? _GEN_111 : writeStack_15_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_400 = alloc ? _GEN_112 : writeStack_16_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_401 = alloc ? _GEN_113 : writeStack_17_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_402 = alloc ? _GEN_114 : writeStack_18_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_403 = alloc ? _GEN_115 : writeStack_19_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_404 = alloc ? _GEN_116 : writeStack_20_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_405 = alloc ? _GEN_117 : writeStack_21_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_406 = alloc ? _GEN_118 : writeStack_22_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_407 = alloc ? _GEN_119 : writeStack_23_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_408 = alloc ? _GEN_120 : writeStack_24_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_409 = alloc ? _GEN_121 : writeStack_25_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_410 = alloc ? _GEN_122 : writeStack_26_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_411 = alloc ? _GEN_123 : writeStack_27_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_412 = alloc ? _GEN_124 : writeStack_28_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_413 = alloc ? _GEN_125 : writeStack_29_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_414 = alloc ? _GEN_126 : writeStack_30_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [1:0] _GEN_415 = alloc ? _GEN_127 : writeStack_31_validStatus; // @[WriteStack.scala 70:14 56:27]
  wire [2:0] _GEN_1856 = {{1'd0}, writeStack_0_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T = _GEN_1856 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_1 = writeStack_0_wvalid & _GEN_1856 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_3 = writeStack_0_wvalid & _GEN_1856 == 3'h1 & writeStack_0_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1857 = {{1'd0}, writeStack_1_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_4 = _GEN_1857 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_5 = writeStack_1_wvalid & _GEN_1857 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_7 = writeStack_1_wvalid & _GEN_1857 == 3'h1 & writeStack_1_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1858 = {{1'd0}, writeStack_2_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_8 = _GEN_1858 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_9 = writeStack_2_wvalid & _GEN_1858 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_11 = writeStack_2_wvalid & _GEN_1858 == 3'h1 & writeStack_2_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1859 = {{1'd0}, writeStack_3_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_12 = _GEN_1859 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_13 = writeStack_3_wvalid & _GEN_1859 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_15 = writeStack_3_wvalid & _GEN_1859 == 3'h1 & writeStack_3_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1860 = {{1'd0}, writeStack_4_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_16 = _GEN_1860 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_17 = writeStack_4_wvalid & _GEN_1860 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_19 = writeStack_4_wvalid & _GEN_1860 == 3'h1 & writeStack_4_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1861 = {{1'd0}, writeStack_5_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_20 = _GEN_1861 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_21 = writeStack_5_wvalid & _GEN_1861 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_23 = writeStack_5_wvalid & _GEN_1861 == 3'h1 & writeStack_5_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1862 = {{1'd0}, writeStack_6_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_24 = _GEN_1862 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_25 = writeStack_6_wvalid & _GEN_1862 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_27 = writeStack_6_wvalid & _GEN_1862 == 3'h1 & writeStack_6_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1863 = {{1'd0}, writeStack_7_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_28 = _GEN_1863 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_29 = writeStack_7_wvalid & _GEN_1863 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_31 = writeStack_7_wvalid & _GEN_1863 == 3'h1 & writeStack_7_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1864 = {{1'd0}, writeStack_8_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_32 = _GEN_1864 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_33 = writeStack_8_wvalid & _GEN_1864 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_35 = writeStack_8_wvalid & _GEN_1864 == 3'h1 & writeStack_8_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1865 = {{1'd0}, writeStack_9_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_36 = _GEN_1865 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_37 = writeStack_9_wvalid & _GEN_1865 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_39 = writeStack_9_wvalid & _GEN_1865 == 3'h1 & writeStack_9_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1866 = {{1'd0}, writeStack_10_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_40 = _GEN_1866 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_41 = writeStack_10_wvalid & _GEN_1866 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_43 = writeStack_10_wvalid & _GEN_1866 == 3'h1 & writeStack_10_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1867 = {{1'd0}, writeStack_11_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_44 = _GEN_1867 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_45 = writeStack_11_wvalid & _GEN_1867 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_47 = writeStack_11_wvalid & _GEN_1867 == 3'h1 & writeStack_11_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1868 = {{1'd0}, writeStack_12_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_48 = _GEN_1868 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_49 = writeStack_12_wvalid & _GEN_1868 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_51 = writeStack_12_wvalid & _GEN_1868 == 3'h1 & writeStack_12_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1869 = {{1'd0}, writeStack_13_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_52 = _GEN_1869 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_53 = writeStack_13_wvalid & _GEN_1869 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_55 = writeStack_13_wvalid & _GEN_1869 == 3'h1 & writeStack_13_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1870 = {{1'd0}, writeStack_14_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_56 = _GEN_1870 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_57 = writeStack_14_wvalid & _GEN_1870 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_59 = writeStack_14_wvalid & _GEN_1870 == 3'h1 & writeStack_14_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1871 = {{1'd0}, writeStack_15_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_60 = _GEN_1871 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_61 = writeStack_15_wvalid & _GEN_1871 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_63 = writeStack_15_wvalid & _GEN_1871 == 3'h1 & writeStack_15_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1872 = {{1'd0}, writeStack_16_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_64 = _GEN_1872 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_65 = writeStack_16_wvalid & _GEN_1872 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_67 = writeStack_16_wvalid & _GEN_1872 == 3'h1 & writeStack_16_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1873 = {{1'd0}, writeStack_17_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_68 = _GEN_1873 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_69 = writeStack_17_wvalid & _GEN_1873 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_71 = writeStack_17_wvalid & _GEN_1873 == 3'h1 & writeStack_17_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1874 = {{1'd0}, writeStack_18_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_72 = _GEN_1874 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_73 = writeStack_18_wvalid & _GEN_1874 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_75 = writeStack_18_wvalid & _GEN_1874 == 3'h1 & writeStack_18_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1875 = {{1'd0}, writeStack_19_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_76 = _GEN_1875 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_77 = writeStack_19_wvalid & _GEN_1875 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_79 = writeStack_19_wvalid & _GEN_1875 == 3'h1 & writeStack_19_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1876 = {{1'd0}, writeStack_20_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_80 = _GEN_1876 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_81 = writeStack_20_wvalid & _GEN_1876 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_83 = writeStack_20_wvalid & _GEN_1876 == 3'h1 & writeStack_20_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1877 = {{1'd0}, writeStack_21_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_84 = _GEN_1877 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_85 = writeStack_21_wvalid & _GEN_1877 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_87 = writeStack_21_wvalid & _GEN_1877 == 3'h1 & writeStack_21_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1878 = {{1'd0}, writeStack_22_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_88 = _GEN_1878 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_89 = writeStack_22_wvalid & _GEN_1878 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_91 = writeStack_22_wvalid & _GEN_1878 == 3'h1 & writeStack_22_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1879 = {{1'd0}, writeStack_23_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_92 = _GEN_1879 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_93 = writeStack_23_wvalid & _GEN_1879 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_95 = writeStack_23_wvalid & _GEN_1879 == 3'h1 & writeStack_23_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1880 = {{1'd0}, writeStack_24_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_96 = _GEN_1880 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_97 = writeStack_24_wvalid & _GEN_1880 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_99 = writeStack_24_wvalid & _GEN_1880 == 3'h1 & writeStack_24_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1881 = {{1'd0}, writeStack_25_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_100 = _GEN_1881 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_101 = writeStack_25_wvalid & _GEN_1881 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_103 = writeStack_25_wvalid & _GEN_1881 == 3'h1 & writeStack_25_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1882 = {{1'd0}, writeStack_26_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_104 = _GEN_1882 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_105 = writeStack_26_wvalid & _GEN_1882 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_107 = writeStack_26_wvalid & _GEN_1882 == 3'h1 & writeStack_26_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1883 = {{1'd0}, writeStack_27_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_108 = _GEN_1883 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_109 = writeStack_27_wvalid & _GEN_1883 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_111 = writeStack_27_wvalid & _GEN_1883 == 3'h1 & writeStack_27_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1884 = {{1'd0}, writeStack_28_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_112 = _GEN_1884 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_113 = writeStack_28_wvalid & _GEN_1884 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_115 = writeStack_28_wvalid & _GEN_1884 == 3'h1 & writeStack_28_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1885 = {{1'd0}, writeStack_29_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_116 = _GEN_1885 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_117 = writeStack_29_wvalid & _GEN_1885 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_119 = writeStack_29_wvalid & _GEN_1885 == 3'h1 & writeStack_29_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1886 = {{1'd0}, writeStack_30_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_120 = _GEN_1886 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_121 = writeStack_30_wvalid & _GEN_1886 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_123 = writeStack_30_wvalid & _GEN_1886 == 3'h1 & writeStack_30_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [2:0] _GEN_1887 = {{1'd0}, writeStack_31_wstatus}; // @[WriteStack.scala 91:60]
  wire  _canW_T_124 = _GEN_1887 == 3'h1; // @[WriteStack.scala 91:60]
  wire  _canW_T_125 = writeStack_31_wvalid & _GEN_1887 == 3'h1; // @[WriteStack.scala 91:47]
  wire  _canW_T_127 = writeStack_31_wvalid & _GEN_1887 == 3'h1 & writeStack_31_waitWFifoId == 5'h0; // @[WriteStack.scala 91:70]
  wire [7:0] canW_lo_lo = {_canW_T_99,_canW_T_103,_canW_T_107,_canW_T_111,_canW_T_115,_canW_T_119,_canW_T_123,
    _canW_T_127}; // @[Cat.scala 31:58]
  wire [15:0] canW_lo = {_canW_T_67,_canW_T_71,_canW_T_75,_canW_T_79,_canW_T_83,_canW_T_87,_canW_T_91,_canW_T_95,
    canW_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] canW_hi_lo = {_canW_T_35,_canW_T_39,_canW_T_43,_canW_T_47,_canW_T_51,_canW_T_55,_canW_T_59,_canW_T_63}; // @[Cat.scala 31:58]
  wire [31:0] _canW_T_128 = {_canW_T_3,_canW_T_7,_canW_T_11,_canW_T_15,_canW_T_19,_canW_T_23,_canW_T_27,_canW_T_31,
    canW_hi_lo,canW_lo}; // @[Cat.scala 31:58]
  wire  _T = io_axiWriteReq_in_aw_ready & io_axiWriteReq_in_aw_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = io_axiWriteReq_in_w_ready & io_axiWriteReq_in_w_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = _T & _T_1; // @[WriteStack.scala 95:34]
  wire [1:0] _writeStack_waitWFifoId_T_64 = _canW_T_1 + _canW_T_5; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_66 = _canW_T_9 + _canW_T_13; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_68 = _writeStack_waitWFifoId_T_64 + _writeStack_waitWFifoId_T_66; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_70 = _canW_T_17 + _canW_T_21; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_72 = _canW_T_25 + _canW_T_29; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_74 = _writeStack_waitWFifoId_T_70 + _writeStack_waitWFifoId_T_72; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_waitWFifoId_T_76 = _writeStack_waitWFifoId_T_68 + _writeStack_waitWFifoId_T_74; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_78 = _canW_T_33 + _canW_T_37; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_80 = _canW_T_41 + _canW_T_45; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_82 = _writeStack_waitWFifoId_T_78 + _writeStack_waitWFifoId_T_80; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_84 = _canW_T_49 + _canW_T_53; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_86 = _canW_T_57 + _canW_T_61; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_88 = _writeStack_waitWFifoId_T_84 + _writeStack_waitWFifoId_T_86; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_waitWFifoId_T_90 = _writeStack_waitWFifoId_T_82 + _writeStack_waitWFifoId_T_88; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_waitWFifoId_T_92 = _writeStack_waitWFifoId_T_76 + _writeStack_waitWFifoId_T_90; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_94 = _canW_T_65 + _canW_T_69; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_96 = _canW_T_73 + _canW_T_77; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_98 = _writeStack_waitWFifoId_T_94 + _writeStack_waitWFifoId_T_96; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_100 = _canW_T_81 + _canW_T_85; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_102 = _canW_T_89 + _canW_T_93; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_104 = _writeStack_waitWFifoId_T_100 + _writeStack_waitWFifoId_T_102; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_waitWFifoId_T_106 = _writeStack_waitWFifoId_T_98 + _writeStack_waitWFifoId_T_104; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_108 = _canW_T_97 + _canW_T_101; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_110 = _canW_T_105 + _canW_T_109; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_112 = _writeStack_waitWFifoId_T_108 + _writeStack_waitWFifoId_T_110; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_114 = _canW_T_113 + _canW_T_117; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_waitWFifoId_T_116 = _canW_T_121 + _canW_T_125; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_waitWFifoId_T_118 = _writeStack_waitWFifoId_T_114 + _writeStack_waitWFifoId_T_116; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_waitWFifoId_T_120 = _writeStack_waitWFifoId_T_112 + _writeStack_waitWFifoId_T_118; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_waitWFifoId_T_122 = _writeStack_waitWFifoId_T_106 + _writeStack_waitWFifoId_T_120; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_waitWFifoId_T_124 = _writeStack_waitWFifoId_T_92 + _writeStack_waitWFifoId_T_122; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_waitWFifoId_T_127 = _writeStack_waitWFifoId_T_124 - 6'h1; // @[WriteStack.scala 98:94]
  wire [4:0] _GEN_576 = 5'h0 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_0_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_577 = 5'h1 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_1_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_578 = 5'h2 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_2_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_579 = 5'h3 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_3_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_580 = 5'h4 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_4_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_581 = 5'h5 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_5_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_582 = 5'h6 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_6_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_583 = 5'h7 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_7_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_584 = 5'h8 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_8_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_585 = 5'h9 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_9_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_586 = 5'ha == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_10_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_587 = 5'hb == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_11_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_588 = 5'hc == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_12_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_589 = 5'hd == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_13_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_590 = 5'he == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_14_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_591 = 5'hf == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_15_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_592 = 5'h10 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_16_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_593 = 5'h11 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_17_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_594 = 5'h12 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_18_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_595 = 5'h13 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_19_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_596 = 5'h14 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_20_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_597 = 5'h15 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_21_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_598 = 5'h16 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_22_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_599 = 5'h17 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_23_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_600 = 5'h18 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_24_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_601 = 5'h19 == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_25_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_602 = 5'h1a == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_26_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_603 = 5'h1b == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_27_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_604 = 5'h1c == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_28_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_605 = 5'h1d == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_29_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_606 = 5'h1e == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_30_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire [4:0] _GEN_607 = 5'h1f == idxInsert ? _writeStack_waitWFifoId_T_127[4:0] : writeStack_31_waitWFifoId; // @[WriteStack.scala 56:27 98:{27,27}]
  wire  _T_6 = _T & ~_T_1; // @[WriteStack.scala 99:44]
  wire [4:0] _GEN_608 = 5'h0 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_0_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_609 = 5'h1 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_1_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_610 = 5'h2 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_2_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_611 = 5'h3 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_3_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_612 = 5'h4 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_4_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_613 = 5'h5 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_5_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_614 = 5'h6 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_6_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_615 = 5'h7 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_7_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_616 = 5'h8 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_8_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_617 = 5'h9 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_9_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_618 = 5'ha == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_10_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_619 = 5'hb == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_11_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_620 = 5'hc == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_12_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_621 = 5'hd == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_13_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_622 = 5'he == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_14_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_623 = 5'hf == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_15_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_624 = 5'h10 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_16_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_625 = 5'h11 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_17_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_626 = 5'h12 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_18_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_627 = 5'h13 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_19_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_628 = 5'h14 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_20_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_629 = 5'h15 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_21_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_630 = 5'h16 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_22_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_631 = 5'h17 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_23_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_632 = 5'h18 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_24_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_633 = 5'h19 == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_25_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_634 = 5'h1a == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_26_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_635 = 5'h1b == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_27_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_636 = 5'h1c == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_28_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_637 = 5'h1d == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_29_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_638 = 5'h1e == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_30_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_639 = 5'h1f == idxInsert ? _writeStack_waitWFifoId_T_124[4:0] : writeStack_31_waitWFifoId; // @[WriteStack.scala 102:{27,27} 56:27]
  wire [4:0] _GEN_640 = _T_6 ? _GEN_608 : writeStack_0_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_641 = _T_6 ? _GEN_609 : writeStack_1_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_642 = _T_6 ? _GEN_610 : writeStack_2_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_643 = _T_6 ? _GEN_611 : writeStack_3_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_644 = _T_6 ? _GEN_612 : writeStack_4_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_645 = _T_6 ? _GEN_613 : writeStack_5_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_646 = _T_6 ? _GEN_614 : writeStack_6_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_647 = _T_6 ? _GEN_615 : writeStack_7_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_648 = _T_6 ? _GEN_616 : writeStack_8_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_649 = _T_6 ? _GEN_617 : writeStack_9_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_650 = _T_6 ? _GEN_618 : writeStack_10_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_651 = _T_6 ? _GEN_619 : writeStack_11_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_652 = _T_6 ? _GEN_620 : writeStack_12_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_653 = _T_6 ? _GEN_621 : writeStack_13_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_654 = _T_6 ? _GEN_622 : writeStack_14_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_655 = _T_6 ? _GEN_623 : writeStack_15_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_656 = _T_6 ? _GEN_624 : writeStack_16_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_657 = _T_6 ? _GEN_625 : writeStack_17_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_658 = _T_6 ? _GEN_626 : writeStack_18_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_659 = _T_6 ? _GEN_627 : writeStack_19_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_660 = _T_6 ? _GEN_628 : writeStack_20_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_661 = _T_6 ? _GEN_629 : writeStack_21_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_662 = _T_6 ? _GEN_630 : writeStack_22_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_663 = _T_6 ? _GEN_631 : writeStack_23_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_664 = _T_6 ? _GEN_632 : writeStack_24_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_665 = _T_6 ? _GEN_633 : writeStack_25_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_666 = _T_6 ? _GEN_634 : writeStack_26_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_667 = _T_6 ? _GEN_635 : writeStack_27_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_668 = _T_6 ? _GEN_636 : writeStack_28_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_669 = _T_6 ? _GEN_637 : writeStack_29_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_670 = _T_6 ? _GEN_638 : writeStack_30_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_671 = _T_6 ? _GEN_639 : writeStack_31_waitWFifoId; // @[WriteStack.scala 100:7 56:27]
  wire [4:0] _GEN_672 = _T_2 ? _GEN_576 : _GEN_640; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_673 = _T_2 ? _GEN_577 : _GEN_641; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_674 = _T_2 ? _GEN_578 : _GEN_642; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_675 = _T_2 ? _GEN_579 : _GEN_643; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_676 = _T_2 ? _GEN_580 : _GEN_644; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_677 = _T_2 ? _GEN_581 : _GEN_645; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_678 = _T_2 ? _GEN_582 : _GEN_646; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_679 = _T_2 ? _GEN_583 : _GEN_647; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_680 = _T_2 ? _GEN_584 : _GEN_648; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_681 = _T_2 ? _GEN_585 : _GEN_649; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_682 = _T_2 ? _GEN_586 : _GEN_650; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_683 = _T_2 ? _GEN_587 : _GEN_651; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_684 = _T_2 ? _GEN_588 : _GEN_652; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_685 = _T_2 ? _GEN_589 : _GEN_653; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_686 = _T_2 ? _GEN_590 : _GEN_654; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_687 = _T_2 ? _GEN_591 : _GEN_655; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_688 = _T_2 ? _GEN_592 : _GEN_656; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_689 = _T_2 ? _GEN_593 : _GEN_657; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_690 = _T_2 ? _GEN_594 : _GEN_658; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_691 = _T_2 ? _GEN_595 : _GEN_659; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_692 = _T_2 ? _GEN_596 : _GEN_660; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_693 = _T_2 ? _GEN_597 : _GEN_661; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_694 = _T_2 ? _GEN_598 : _GEN_662; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_695 = _T_2 ? _GEN_599 : _GEN_663; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_696 = _T_2 ? _GEN_600 : _GEN_664; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_697 = _T_2 ? _GEN_601 : _GEN_665; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_698 = _T_2 ? _GEN_602 : _GEN_666; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_699 = _T_2 ? _GEN_603 : _GEN_667; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_700 = _T_2 ? _GEN_604 : _GEN_668; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_701 = _T_2 ? _GEN_605 : _GEN_669; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_702 = _T_2 ? _GEN_606 : _GEN_670; // @[WriteStack.scala 96:7]
  wire [4:0] _GEN_703 = _T_2 ? _GEN_607 : _GEN_671; // @[WriteStack.scala 96:7]
  wire [4:0] _writeStack_0_waitWFifoId_T_1 = writeStack_0_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_707 = _canW_T_3 ? 3'h2 : {{1'd0}, _GEN_352}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_1_waitWFifoId_T_1 = writeStack_1_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_712 = _canW_T_7 ? 3'h2 : {{1'd0}, _GEN_353}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_2_waitWFifoId_T_1 = writeStack_2_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_717 = _canW_T_11 ? 3'h2 : {{1'd0}, _GEN_354}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_3_waitWFifoId_T_1 = writeStack_3_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_722 = _canW_T_15 ? 3'h2 : {{1'd0}, _GEN_355}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_4_waitWFifoId_T_1 = writeStack_4_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_727 = _canW_T_19 ? 3'h2 : {{1'd0}, _GEN_356}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_5_waitWFifoId_T_1 = writeStack_5_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_732 = _canW_T_23 ? 3'h2 : {{1'd0}, _GEN_357}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_6_waitWFifoId_T_1 = writeStack_6_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_737 = _canW_T_27 ? 3'h2 : {{1'd0}, _GEN_358}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_7_waitWFifoId_T_1 = writeStack_7_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_742 = _canW_T_31 ? 3'h2 : {{1'd0}, _GEN_359}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_8_waitWFifoId_T_1 = writeStack_8_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_747 = _canW_T_35 ? 3'h2 : {{1'd0}, _GEN_360}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_9_waitWFifoId_T_1 = writeStack_9_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_752 = _canW_T_39 ? 3'h2 : {{1'd0}, _GEN_361}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_10_waitWFifoId_T_1 = writeStack_10_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_757 = _canW_T_43 ? 3'h2 : {{1'd0}, _GEN_362}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_11_waitWFifoId_T_1 = writeStack_11_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_762 = _canW_T_47 ? 3'h2 : {{1'd0}, _GEN_363}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_12_waitWFifoId_T_1 = writeStack_12_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_767 = _canW_T_51 ? 3'h2 : {{1'd0}, _GEN_364}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_13_waitWFifoId_T_1 = writeStack_13_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_772 = _canW_T_55 ? 3'h2 : {{1'd0}, _GEN_365}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_14_waitWFifoId_T_1 = writeStack_14_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_777 = _canW_T_59 ? 3'h2 : {{1'd0}, _GEN_366}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_15_waitWFifoId_T_1 = writeStack_15_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_782 = _canW_T_63 ? 3'h2 : {{1'd0}, _GEN_367}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_16_waitWFifoId_T_1 = writeStack_16_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_787 = _canW_T_67 ? 3'h2 : {{1'd0}, _GEN_368}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_17_waitWFifoId_T_1 = writeStack_17_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_792 = _canW_T_71 ? 3'h2 : {{1'd0}, _GEN_369}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_18_waitWFifoId_T_1 = writeStack_18_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_797 = _canW_T_75 ? 3'h2 : {{1'd0}, _GEN_370}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_19_waitWFifoId_T_1 = writeStack_19_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_802 = _canW_T_79 ? 3'h2 : {{1'd0}, _GEN_371}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_20_waitWFifoId_T_1 = writeStack_20_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_807 = _canW_T_83 ? 3'h2 : {{1'd0}, _GEN_372}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_21_waitWFifoId_T_1 = writeStack_21_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_812 = _canW_T_87 ? 3'h2 : {{1'd0}, _GEN_373}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_22_waitWFifoId_T_1 = writeStack_22_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_817 = _canW_T_91 ? 3'h2 : {{1'd0}, _GEN_374}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_23_waitWFifoId_T_1 = writeStack_23_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_822 = _canW_T_95 ? 3'h2 : {{1'd0}, _GEN_375}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_24_waitWFifoId_T_1 = writeStack_24_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_827 = _canW_T_99 ? 3'h2 : {{1'd0}, _GEN_376}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_25_waitWFifoId_T_1 = writeStack_25_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_832 = _canW_T_103 ? 3'h2 : {{1'd0}, _GEN_377}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_26_waitWFifoId_T_1 = writeStack_26_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_837 = _canW_T_107 ? 3'h2 : {{1'd0}, _GEN_378}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_27_waitWFifoId_T_1 = writeStack_27_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_842 = _canW_T_111 ? 3'h2 : {{1'd0}, _GEN_379}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_28_waitWFifoId_T_1 = writeStack_28_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_847 = _canW_T_115 ? 3'h2 : {{1'd0}, _GEN_380}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_29_waitWFifoId_T_1 = writeStack_29_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_852 = _canW_T_119 ? 3'h2 : {{1'd0}, _GEN_381}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_30_waitWFifoId_T_1 = writeStack_30_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_857 = _canW_T_123 ? 3'h2 : {{1'd0}, _GEN_382}; // @[WriteStack.scala 109:76 112:27]
  wire [4:0] _writeStack_31_waitWFifoId_T_1 = writeStack_31_waitWFifoId - 5'h1; // @[WriteStack.scala 113:47]
  wire [2:0] _GEN_862 = _canW_T_127 ? 3'h2 : {{1'd0}, _GEN_383}; // @[WriteStack.scala 109:76 112:27]
  wire [2:0] _GEN_866 = _T_1 ? _GEN_707 : {{1'd0}, _GEN_352}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_870 = _T_1 ? _GEN_712 : {{1'd0}, _GEN_353}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_874 = _T_1 ? _GEN_717 : {{1'd0}, _GEN_354}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_878 = _T_1 ? _GEN_722 : {{1'd0}, _GEN_355}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_882 = _T_1 ? _GEN_727 : {{1'd0}, _GEN_356}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_886 = _T_1 ? _GEN_732 : {{1'd0}, _GEN_357}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_890 = _T_1 ? _GEN_737 : {{1'd0}, _GEN_358}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_894 = _T_1 ? _GEN_742 : {{1'd0}, _GEN_359}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_898 = _T_1 ? _GEN_747 : {{1'd0}, _GEN_360}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_902 = _T_1 ? _GEN_752 : {{1'd0}, _GEN_361}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_906 = _T_1 ? _GEN_757 : {{1'd0}, _GEN_362}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_910 = _T_1 ? _GEN_762 : {{1'd0}, _GEN_363}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_914 = _T_1 ? _GEN_767 : {{1'd0}, _GEN_364}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_918 = _T_1 ? _GEN_772 : {{1'd0}, _GEN_365}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_922 = _T_1 ? _GEN_777 : {{1'd0}, _GEN_366}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_926 = _T_1 ? _GEN_782 : {{1'd0}, _GEN_367}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_930 = _T_1 ? _GEN_787 : {{1'd0}, _GEN_368}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_934 = _T_1 ? _GEN_792 : {{1'd0}, _GEN_369}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_938 = _T_1 ? _GEN_797 : {{1'd0}, _GEN_370}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_942 = _T_1 ? _GEN_802 : {{1'd0}, _GEN_371}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_946 = _T_1 ? _GEN_807 : {{1'd0}, _GEN_372}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_950 = _T_1 ? _GEN_812 : {{1'd0}, _GEN_373}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_954 = _T_1 ? _GEN_817 : {{1'd0}, _GEN_374}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_958 = _T_1 ? _GEN_822 : {{1'd0}, _GEN_375}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_962 = _T_1 ? _GEN_827 : {{1'd0}, _GEN_376}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_966 = _T_1 ? _GEN_832 : {{1'd0}, _GEN_377}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_970 = _T_1 ? _GEN_837 : {{1'd0}, _GEN_378}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_974 = _T_1 ? _GEN_842 : {{1'd0}, _GEN_379}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_978 = _T_1 ? _GEN_847 : {{1'd0}, _GEN_380}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_982 = _T_1 ? _GEN_852 : {{1'd0}, _GEN_381}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_986 = _T_1 ? _GEN_857 : {{1'd0}, _GEN_382}; // @[WriteStack.scala 106:5]
  wire [2:0] _GEN_990 = _T_1 ? _GEN_862 : {{1'd0}, _GEN_383}; // @[WriteStack.scala 106:5]
  wire  _hasValid_T = writeStack_0_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_1 = writeStack_0_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_2 = writeStack_0_validStatus == 2'h1 & writeStack_0_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_3 = writeStack_1_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_4 = writeStack_1_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_5 = writeStack_1_validStatus == 2'h1 & writeStack_1_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_6 = writeStack_2_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_7 = writeStack_2_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_8 = writeStack_2_validStatus == 2'h1 & writeStack_2_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_9 = writeStack_3_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_10 = writeStack_3_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_11 = writeStack_3_validStatus == 2'h1 & writeStack_3_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_12 = writeStack_4_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_13 = writeStack_4_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_14 = writeStack_4_validStatus == 2'h1 & writeStack_4_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_15 = writeStack_5_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_16 = writeStack_5_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_17 = writeStack_5_validStatus == 2'h1 & writeStack_5_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_18 = writeStack_6_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_19 = writeStack_6_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_20 = writeStack_6_validStatus == 2'h1 & writeStack_6_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_21 = writeStack_7_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_22 = writeStack_7_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_23 = writeStack_7_validStatus == 2'h1 & writeStack_7_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_24 = writeStack_8_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_25 = writeStack_8_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_26 = writeStack_8_validStatus == 2'h1 & writeStack_8_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_27 = writeStack_9_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_28 = writeStack_9_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_29 = writeStack_9_validStatus == 2'h1 & writeStack_9_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_30 = writeStack_10_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_31 = writeStack_10_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_32 = writeStack_10_validStatus == 2'h1 & writeStack_10_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_33 = writeStack_11_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_34 = writeStack_11_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_35 = writeStack_11_validStatus == 2'h1 & writeStack_11_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_36 = writeStack_12_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_37 = writeStack_12_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_38 = writeStack_12_validStatus == 2'h1 & writeStack_12_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_39 = writeStack_13_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_40 = writeStack_13_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_41 = writeStack_13_validStatus == 2'h1 & writeStack_13_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_42 = writeStack_14_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_43 = writeStack_14_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_44 = writeStack_14_validStatus == 2'h1 & writeStack_14_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_45 = writeStack_15_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_46 = writeStack_15_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_47 = writeStack_15_validStatus == 2'h1 & writeStack_15_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_48 = writeStack_16_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_49 = writeStack_16_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_50 = writeStack_16_validStatus == 2'h1 & writeStack_16_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_51 = writeStack_17_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_52 = writeStack_17_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_53 = writeStack_17_validStatus == 2'h1 & writeStack_17_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_54 = writeStack_18_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_55 = writeStack_18_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_56 = writeStack_18_validStatus == 2'h1 & writeStack_18_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_57 = writeStack_19_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_58 = writeStack_19_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_59 = writeStack_19_validStatus == 2'h1 & writeStack_19_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_60 = writeStack_20_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_61 = writeStack_20_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_62 = writeStack_20_validStatus == 2'h1 & writeStack_20_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_63 = writeStack_21_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_64 = writeStack_21_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_65 = writeStack_21_validStatus == 2'h1 & writeStack_21_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_66 = writeStack_22_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_67 = writeStack_22_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_68 = writeStack_22_validStatus == 2'h1 & writeStack_22_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_69 = writeStack_23_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_70 = writeStack_23_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_71 = writeStack_23_validStatus == 2'h1 & writeStack_23_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_72 = writeStack_24_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_73 = writeStack_24_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_74 = writeStack_24_validStatus == 2'h1 & writeStack_24_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_75 = writeStack_25_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_76 = writeStack_25_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_77 = writeStack_25_validStatus == 2'h1 & writeStack_25_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_78 = writeStack_26_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_79 = writeStack_26_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_80 = writeStack_26_validStatus == 2'h1 & writeStack_26_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_81 = writeStack_27_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_82 = writeStack_27_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_83 = writeStack_27_validStatus == 2'h1 & writeStack_27_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_84 = writeStack_28_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_85 = writeStack_28_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_86 = writeStack_28_validStatus == 2'h1 & writeStack_28_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_87 = writeStack_29_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_88 = writeStack_29_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_89 = writeStack_29_validStatus == 2'h1 & writeStack_29_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_90 = writeStack_30_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_91 = writeStack_30_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_92 = writeStack_30_validStatus == 2'h1 & writeStack_30_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _hasValid_T_93 = writeStack_31_validStatus == 2'h1; // @[WriteStack.scala 122:57]
  wire  _hasValid_T_94 = writeStack_31_validFifoId == 5'h0; // @[WriteStack.scala 122:88]
  wire  _hasValid_T_95 = writeStack_31_validStatus == 2'h1 & writeStack_31_validFifoId == 5'h0; // @[WriteStack.scala 122:71]
  wire  _T_201 = io_validReq_in_ready & io_validReq_in_valid; // @[Decoupled.scala 50:35]
  wire  _T_202 = _T & _T_201; // @[WriteStack.scala 138:34]
  wire  _writeStack_validFifoId_T_1 = writeStack_0_wvalid & _hasValid_T; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_3 = writeStack_1_wvalid & _hasValid_T_3; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_5 = writeStack_2_wvalid & _hasValid_T_6; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_7 = writeStack_3_wvalid & _hasValid_T_9; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_9 = writeStack_4_wvalid & _hasValid_T_12; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_11 = writeStack_5_wvalid & _hasValid_T_15; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_13 = writeStack_6_wvalid & _hasValid_T_18; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_15 = writeStack_7_wvalid & _hasValid_T_21; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_17 = writeStack_8_wvalid & _hasValid_T_24; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_19 = writeStack_9_wvalid & _hasValid_T_27; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_21 = writeStack_10_wvalid & _hasValid_T_30; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_23 = writeStack_11_wvalid & _hasValid_T_33; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_25 = writeStack_12_wvalid & _hasValid_T_36; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_27 = writeStack_13_wvalid & _hasValid_T_39; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_29 = writeStack_14_wvalid & _hasValid_T_42; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_31 = writeStack_15_wvalid & _hasValid_T_45; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_33 = writeStack_16_wvalid & _hasValid_T_48; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_35 = writeStack_17_wvalid & _hasValid_T_51; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_37 = writeStack_18_wvalid & _hasValid_T_54; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_39 = writeStack_19_wvalid & _hasValid_T_57; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_41 = writeStack_20_wvalid & _hasValid_T_60; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_43 = writeStack_21_wvalid & _hasValid_T_63; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_45 = writeStack_22_wvalid & _hasValid_T_66; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_47 = writeStack_23_wvalid & _hasValid_T_69; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_49 = writeStack_24_wvalid & _hasValid_T_72; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_51 = writeStack_25_wvalid & _hasValid_T_75; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_53 = writeStack_26_wvalid & _hasValid_T_78; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_55 = writeStack_27_wvalid & _hasValid_T_81; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_57 = writeStack_28_wvalid & _hasValid_T_84; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_59 = writeStack_29_wvalid & _hasValid_T_87; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_61 = writeStack_30_wvalid & _hasValid_T_90; // @[WriteStack.scala 141:67]
  wire  _writeStack_validFifoId_T_63 = writeStack_31_wvalid & _hasValid_T_93; // @[WriteStack.scala 141:67]
  wire [1:0] _writeStack_validFifoId_T_64 = _writeStack_validFifoId_T_1 + _writeStack_validFifoId_T_3; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_66 = _writeStack_validFifoId_T_5 + _writeStack_validFifoId_T_7; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_68 = _writeStack_validFifoId_T_64 + _writeStack_validFifoId_T_66; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_70 = _writeStack_validFifoId_T_9 + _writeStack_validFifoId_T_11; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_72 = _writeStack_validFifoId_T_13 + _writeStack_validFifoId_T_15; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_74 = _writeStack_validFifoId_T_70 + _writeStack_validFifoId_T_72; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_validFifoId_T_76 = _writeStack_validFifoId_T_68 + _writeStack_validFifoId_T_74; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_78 = _writeStack_validFifoId_T_17 + _writeStack_validFifoId_T_19; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_80 = _writeStack_validFifoId_T_21 + _writeStack_validFifoId_T_23; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_82 = _writeStack_validFifoId_T_78 + _writeStack_validFifoId_T_80; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_84 = _writeStack_validFifoId_T_25 + _writeStack_validFifoId_T_27; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_86 = _writeStack_validFifoId_T_29 + _writeStack_validFifoId_T_31; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_88 = _writeStack_validFifoId_T_84 + _writeStack_validFifoId_T_86; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_validFifoId_T_90 = _writeStack_validFifoId_T_82 + _writeStack_validFifoId_T_88; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_validFifoId_T_92 = _writeStack_validFifoId_T_76 + _writeStack_validFifoId_T_90; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_94 = _writeStack_validFifoId_T_33 + _writeStack_validFifoId_T_35; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_96 = _writeStack_validFifoId_T_37 + _writeStack_validFifoId_T_39; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_98 = _writeStack_validFifoId_T_94 + _writeStack_validFifoId_T_96; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_100 = _writeStack_validFifoId_T_41 + _writeStack_validFifoId_T_43; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_102 = _writeStack_validFifoId_T_45 + _writeStack_validFifoId_T_47; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_104 = _writeStack_validFifoId_T_100 + _writeStack_validFifoId_T_102; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_validFifoId_T_106 = _writeStack_validFifoId_T_98 + _writeStack_validFifoId_T_104; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_108 = _writeStack_validFifoId_T_49 + _writeStack_validFifoId_T_51; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_110 = _writeStack_validFifoId_T_53 + _writeStack_validFifoId_T_55; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_112 = _writeStack_validFifoId_T_108 + _writeStack_validFifoId_T_110; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_114 = _writeStack_validFifoId_T_57 + _writeStack_validFifoId_T_59; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_validFifoId_T_116 = _writeStack_validFifoId_T_61 + _writeStack_validFifoId_T_63; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_validFifoId_T_118 = _writeStack_validFifoId_T_114 + _writeStack_validFifoId_T_116; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_validFifoId_T_120 = _writeStack_validFifoId_T_112 + _writeStack_validFifoId_T_118; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_validFifoId_T_122 = _writeStack_validFifoId_T_106 + _writeStack_validFifoId_T_120; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_validFifoId_T_124 = _writeStack_validFifoId_T_92 + _writeStack_validFifoId_T_122; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_validFifoId_T_127 = _writeStack_validFifoId_T_124 - 6'h1; // @[WriteStack.scala 141:102]
  wire [4:0] _GEN_992 = 5'h0 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_0_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_993 = 5'h1 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_1_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_994 = 5'h2 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_2_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_995 = 5'h3 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_3_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_996 = 5'h4 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_4_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_997 = 5'h5 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_5_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_998 = 5'h6 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_6_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_999 = 5'h7 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_7_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1000 = 5'h8 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_8_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1001 = 5'h9 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_9_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1002 = 5'ha == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_10_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1003 = 5'hb == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_11_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1004 = 5'hc == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_12_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1005 = 5'hd == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_13_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1006 = 5'he == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_14_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1007 = 5'hf == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_15_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1008 = 5'h10 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_16_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1009 = 5'h11 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_17_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1010 = 5'h12 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_18_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1011 = 5'h13 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_19_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1012 = 5'h14 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_20_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1013 = 5'h15 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_21_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1014 = 5'h16 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_22_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1015 = 5'h17 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_23_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1016 = 5'h18 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_24_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1017 = 5'h19 == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_25_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1018 = 5'h1a == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_26_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1019 = 5'h1b == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_27_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1020 = 5'h1c == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_28_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1021 = 5'h1d == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_29_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1022 = 5'h1e == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_30_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire [4:0] _GEN_1023 = 5'h1f == idxInsert ? _writeStack_validFifoId_T_127[4:0] : writeStack_31_validFifoId; // @[WriteStack.scala 141:{27,27} 56:27]
  wire  _T_206 = _T & ~_T_201; // @[WriteStack.scala 142:44]
  wire [4:0] _GEN_1024 = 5'h0 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_0_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1025 = 5'h1 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_1_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1026 = 5'h2 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_2_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1027 = 5'h3 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_3_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1028 = 5'h4 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_4_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1029 = 5'h5 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_5_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1030 = 5'h6 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_6_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1031 = 5'h7 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_7_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1032 = 5'h8 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_8_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1033 = 5'h9 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_9_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1034 = 5'ha == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_10_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1035 = 5'hb == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_11_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1036 = 5'hc == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_12_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1037 = 5'hd == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_13_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1038 = 5'he == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_14_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1039 = 5'hf == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_15_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1040 = 5'h10 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_16_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1041 = 5'h11 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_17_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1042 = 5'h12 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_18_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1043 = 5'h13 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_19_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1044 = 5'h14 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_20_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1045 = 5'h15 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_21_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1046 = 5'h16 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_22_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1047 = 5'h17 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_23_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1048 = 5'h18 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_24_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1049 = 5'h19 == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_25_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1050 = 5'h1a == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_26_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1051 = 5'h1b == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_27_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1052 = 5'h1c == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_28_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1053 = 5'h1d == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_29_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1054 = 5'h1e == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_30_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1055 = 5'h1f == idxInsert ? _writeStack_validFifoId_T_124[4:0] : writeStack_31_validFifoId; // @[WriteStack.scala 145:{27,27} 56:27]
  wire [4:0] _GEN_1056 = _T_206 ? _GEN_1024 : writeStack_0_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1057 = _T_206 ? _GEN_1025 : writeStack_1_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1058 = _T_206 ? _GEN_1026 : writeStack_2_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1059 = _T_206 ? _GEN_1027 : writeStack_3_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1060 = _T_206 ? _GEN_1028 : writeStack_4_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1061 = _T_206 ? _GEN_1029 : writeStack_5_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1062 = _T_206 ? _GEN_1030 : writeStack_6_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1063 = _T_206 ? _GEN_1031 : writeStack_7_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1064 = _T_206 ? _GEN_1032 : writeStack_8_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1065 = _T_206 ? _GEN_1033 : writeStack_9_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1066 = _T_206 ? _GEN_1034 : writeStack_10_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1067 = _T_206 ? _GEN_1035 : writeStack_11_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1068 = _T_206 ? _GEN_1036 : writeStack_12_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1069 = _T_206 ? _GEN_1037 : writeStack_13_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1070 = _T_206 ? _GEN_1038 : writeStack_14_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1071 = _T_206 ? _GEN_1039 : writeStack_15_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1072 = _T_206 ? _GEN_1040 : writeStack_16_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1073 = _T_206 ? _GEN_1041 : writeStack_17_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1074 = _T_206 ? _GEN_1042 : writeStack_18_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1075 = _T_206 ? _GEN_1043 : writeStack_19_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1076 = _T_206 ? _GEN_1044 : writeStack_20_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1077 = _T_206 ? _GEN_1045 : writeStack_21_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1078 = _T_206 ? _GEN_1046 : writeStack_22_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1079 = _T_206 ? _GEN_1047 : writeStack_23_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1080 = _T_206 ? _GEN_1048 : writeStack_24_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1081 = _T_206 ? _GEN_1049 : writeStack_25_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1082 = _T_206 ? _GEN_1050 : writeStack_26_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1083 = _T_206 ? _GEN_1051 : writeStack_27_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1084 = _T_206 ? _GEN_1052 : writeStack_28_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1085 = _T_206 ? _GEN_1053 : writeStack_29_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1086 = _T_206 ? _GEN_1054 : writeStack_30_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1087 = _T_206 ? _GEN_1055 : writeStack_31_validFifoId; // @[WriteStack.scala 143:7 56:27]
  wire [4:0] _GEN_1088 = _T_202 ? _GEN_992 : _GEN_1056; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1089 = _T_202 ? _GEN_993 : _GEN_1057; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1090 = _T_202 ? _GEN_994 : _GEN_1058; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1091 = _T_202 ? _GEN_995 : _GEN_1059; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1092 = _T_202 ? _GEN_996 : _GEN_1060; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1093 = _T_202 ? _GEN_997 : _GEN_1061; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1094 = _T_202 ? _GEN_998 : _GEN_1062; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1095 = _T_202 ? _GEN_999 : _GEN_1063; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1096 = _T_202 ? _GEN_1000 : _GEN_1064; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1097 = _T_202 ? _GEN_1001 : _GEN_1065; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1098 = _T_202 ? _GEN_1002 : _GEN_1066; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1099 = _T_202 ? _GEN_1003 : _GEN_1067; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1100 = _T_202 ? _GEN_1004 : _GEN_1068; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1101 = _T_202 ? _GEN_1005 : _GEN_1069; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1102 = _T_202 ? _GEN_1006 : _GEN_1070; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1103 = _T_202 ? _GEN_1007 : _GEN_1071; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1104 = _T_202 ? _GEN_1008 : _GEN_1072; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1105 = _T_202 ? _GEN_1009 : _GEN_1073; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1106 = _T_202 ? _GEN_1010 : _GEN_1074; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1107 = _T_202 ? _GEN_1011 : _GEN_1075; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1108 = _T_202 ? _GEN_1012 : _GEN_1076; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1109 = _T_202 ? _GEN_1013 : _GEN_1077; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1110 = _T_202 ? _GEN_1014 : _GEN_1078; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1111 = _T_202 ? _GEN_1015 : _GEN_1079; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1112 = _T_202 ? _GEN_1016 : _GEN_1080; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1113 = _T_202 ? _GEN_1017 : _GEN_1081; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1114 = _T_202 ? _GEN_1018 : _GEN_1082; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1115 = _T_202 ? _GEN_1019 : _GEN_1083; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1116 = _T_202 ? _GEN_1020 : _GEN_1084; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1117 = _T_202 ? _GEN_1021 : _GEN_1085; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1118 = _T_202 ? _GEN_1022 : _GEN_1086; // @[WriteStack.scala 139:7]
  wire [4:0] _GEN_1119 = _T_202 ? _GEN_1023 : _GEN_1087; // @[WriteStack.scala 139:7]
  wire [4:0] _writeStack_0_validFifoId_T_1 = writeStack_0_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1121 = _writeStack_validFifoId_T_1 & _hasValid_T_1 ? 2'h2 : _GEN_384; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_1_validFifoId_T_1 = writeStack_1_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1124 = _writeStack_validFifoId_T_3 & _hasValid_T_4 ? 2'h2 : _GEN_385; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_2_validFifoId_T_1 = writeStack_2_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1127 = _writeStack_validFifoId_T_5 & _hasValid_T_7 ? 2'h2 : _GEN_386; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_3_validFifoId_T_1 = writeStack_3_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1130 = _writeStack_validFifoId_T_7 & _hasValid_T_10 ? 2'h2 : _GEN_387; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_4_validFifoId_T_1 = writeStack_4_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1133 = _writeStack_validFifoId_T_9 & _hasValid_T_13 ? 2'h2 : _GEN_388; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_5_validFifoId_T_1 = writeStack_5_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1136 = _writeStack_validFifoId_T_11 & _hasValid_T_16 ? 2'h2 : _GEN_389; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_6_validFifoId_T_1 = writeStack_6_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1139 = _writeStack_validFifoId_T_13 & _hasValid_T_19 ? 2'h2 : _GEN_390; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_7_validFifoId_T_1 = writeStack_7_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1142 = _writeStack_validFifoId_T_15 & _hasValid_T_22 ? 2'h2 : _GEN_391; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_8_validFifoId_T_1 = writeStack_8_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1145 = _writeStack_validFifoId_T_17 & _hasValid_T_25 ? 2'h2 : _GEN_392; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_9_validFifoId_T_1 = writeStack_9_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1148 = _writeStack_validFifoId_T_19 & _hasValid_T_28 ? 2'h2 : _GEN_393; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_10_validFifoId_T_1 = writeStack_10_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1151 = _writeStack_validFifoId_T_21 & _hasValid_T_31 ? 2'h2 : _GEN_394; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_11_validFifoId_T_1 = writeStack_11_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1154 = _writeStack_validFifoId_T_23 & _hasValid_T_34 ? 2'h2 : _GEN_395; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_12_validFifoId_T_1 = writeStack_12_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1157 = _writeStack_validFifoId_T_25 & _hasValid_T_37 ? 2'h2 : _GEN_396; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_13_validFifoId_T_1 = writeStack_13_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1160 = _writeStack_validFifoId_T_27 & _hasValid_T_40 ? 2'h2 : _GEN_397; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_14_validFifoId_T_1 = writeStack_14_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1163 = _writeStack_validFifoId_T_29 & _hasValid_T_43 ? 2'h2 : _GEN_398; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_15_validFifoId_T_1 = writeStack_15_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1166 = _writeStack_validFifoId_T_31 & _hasValid_T_46 ? 2'h2 : _GEN_399; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_16_validFifoId_T_1 = writeStack_16_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1169 = _writeStack_validFifoId_T_33 & _hasValid_T_49 ? 2'h2 : _GEN_400; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_17_validFifoId_T_1 = writeStack_17_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1172 = _writeStack_validFifoId_T_35 & _hasValid_T_52 ? 2'h2 : _GEN_401; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_18_validFifoId_T_1 = writeStack_18_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1175 = _writeStack_validFifoId_T_37 & _hasValid_T_55 ? 2'h2 : _GEN_402; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_19_validFifoId_T_1 = writeStack_19_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1178 = _writeStack_validFifoId_T_39 & _hasValid_T_58 ? 2'h2 : _GEN_403; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_20_validFifoId_T_1 = writeStack_20_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1181 = _writeStack_validFifoId_T_41 & _hasValid_T_61 ? 2'h2 : _GEN_404; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_21_validFifoId_T_1 = writeStack_21_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1184 = _writeStack_validFifoId_T_43 & _hasValid_T_64 ? 2'h2 : _GEN_405; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_22_validFifoId_T_1 = writeStack_22_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1187 = _writeStack_validFifoId_T_45 & _hasValid_T_67 ? 2'h2 : _GEN_406; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_23_validFifoId_T_1 = writeStack_23_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1190 = _writeStack_validFifoId_T_47 & _hasValid_T_70 ? 2'h2 : _GEN_407; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_24_validFifoId_T_1 = writeStack_24_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1193 = _writeStack_validFifoId_T_49 & _hasValid_T_73 ? 2'h2 : _GEN_408; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_25_validFifoId_T_1 = writeStack_25_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1196 = _writeStack_validFifoId_T_51 & _hasValid_T_76 ? 2'h2 : _GEN_409; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_26_validFifoId_T_1 = writeStack_26_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1199 = _writeStack_validFifoId_T_53 & _hasValid_T_79 ? 2'h2 : _GEN_410; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_27_validFifoId_T_1 = writeStack_27_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1202 = _writeStack_validFifoId_T_55 & _hasValid_T_82 ? 2'h2 : _GEN_411; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_28_validFifoId_T_1 = writeStack_28_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1205 = _writeStack_validFifoId_T_57 & _hasValid_T_85 ? 2'h2 : _GEN_412; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_29_validFifoId_T_1 = writeStack_29_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1208 = _writeStack_validFifoId_T_59 & _hasValid_T_88 ? 2'h2 : _GEN_413; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_30_validFifoId_T_1 = writeStack_30_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1211 = _writeStack_validFifoId_T_61 & _hasValid_T_91 ? 2'h2 : _GEN_414; // @[WriteStack.scala 151:84 152:29]
  wire [4:0] _writeStack_31_validFifoId_T_1 = writeStack_31_validFifoId - 5'h1; // @[WriteStack.scala 153:46]
  wire [1:0] _GEN_1214 = _writeStack_validFifoId_T_63 & _hasValid_T_94 ? 2'h2 : _GEN_415; // @[WriteStack.scala 151:84 152:29]
  wire [1:0] _GEN_1216 = _T_201 ? _GEN_1121 : _GEN_384; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1218 = _T_201 ? _GEN_1124 : _GEN_385; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1220 = _T_201 ? _GEN_1127 : _GEN_386; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1222 = _T_201 ? _GEN_1130 : _GEN_387; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1224 = _T_201 ? _GEN_1133 : _GEN_388; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1226 = _T_201 ? _GEN_1136 : _GEN_389; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1228 = _T_201 ? _GEN_1139 : _GEN_390; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1230 = _T_201 ? _GEN_1142 : _GEN_391; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1232 = _T_201 ? _GEN_1145 : _GEN_392; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1234 = _T_201 ? _GEN_1148 : _GEN_393; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1236 = _T_201 ? _GEN_1151 : _GEN_394; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1238 = _T_201 ? _GEN_1154 : _GEN_395; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1240 = _T_201 ? _GEN_1157 : _GEN_396; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1242 = _T_201 ? _GEN_1160 : _GEN_397; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1244 = _T_201 ? _GEN_1163 : _GEN_398; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1246 = _T_201 ? _GEN_1166 : _GEN_399; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1248 = _T_201 ? _GEN_1169 : _GEN_400; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1250 = _T_201 ? _GEN_1172 : _GEN_401; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1252 = _T_201 ? _GEN_1175 : _GEN_402; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1254 = _T_201 ? _GEN_1178 : _GEN_403; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1256 = _T_201 ? _GEN_1181 : _GEN_404; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1258 = _T_201 ? _GEN_1184 : _GEN_405; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1260 = _T_201 ? _GEN_1187 : _GEN_406; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1262 = _T_201 ? _GEN_1190 : _GEN_407; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1264 = _T_201 ? _GEN_1193 : _GEN_408; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1266 = _T_201 ? _GEN_1196 : _GEN_409; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1268 = _T_201 ? _GEN_1199 : _GEN_410; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1270 = _T_201 ? _GEN_1202 : _GEN_411; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1272 = _T_201 ? _GEN_1205 : _GEN_412; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1274 = _T_201 ? _GEN_1208 : _GEN_413; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1276 = _T_201 ? _GEN_1211 : _GEN_414; // @[WriteStack.scala 148:5]
  wire [1:0] _GEN_1278 = _T_201 ? _GEN_1214 : _GEN_415; // @[WriteStack.scala 148:5]
  wire  _canValid_T_1 = writeStack_0_wvalid & writeStack_0_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_3 = writeStack_1_wvalid & writeStack_1_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_5 = writeStack_2_wvalid & writeStack_2_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_7 = writeStack_3_wvalid & writeStack_3_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_9 = writeStack_4_wvalid & writeStack_4_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_11 = writeStack_5_wvalid & writeStack_5_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_13 = writeStack_6_wvalid & writeStack_6_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_15 = writeStack_7_wvalid & writeStack_7_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_17 = writeStack_8_wvalid & writeStack_8_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_19 = writeStack_9_wvalid & writeStack_9_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_21 = writeStack_10_wvalid & writeStack_10_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_23 = writeStack_11_wvalid & writeStack_11_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_25 = writeStack_12_wvalid & writeStack_12_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_27 = writeStack_13_wvalid & writeStack_13_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_29 = writeStack_14_wvalid & writeStack_14_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_31 = writeStack_15_wvalid & writeStack_15_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_33 = writeStack_16_wvalid & writeStack_16_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_35 = writeStack_17_wvalid & writeStack_17_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_37 = writeStack_18_wvalid & writeStack_18_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_39 = writeStack_19_wvalid & writeStack_19_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_41 = writeStack_20_wvalid & writeStack_20_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_43 = writeStack_21_wvalid & writeStack_21_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_45 = writeStack_22_wvalid & writeStack_22_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_47 = writeStack_23_wvalid & writeStack_23_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_49 = writeStack_24_wvalid & writeStack_24_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_51 = writeStack_25_wvalid & writeStack_25_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_53 = writeStack_26_wvalid & writeStack_26_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_55 = writeStack_27_wvalid & writeStack_27_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_57 = writeStack_28_wvalid & writeStack_28_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_59 = writeStack_29_wvalid & writeStack_29_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_61 = writeStack_30_wvalid & writeStack_30_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire  _canValid_T_63 = writeStack_31_wvalid & writeStack_31_validStatus == 2'h2; // @[WriteStack.scala 162:51]
  wire [7:0] canValid_lo_lo = {_canValid_T_49,_canValid_T_51,_canValid_T_53,_canValid_T_55,_canValid_T_57,_canValid_T_59
    ,_canValid_T_61,_canValid_T_63}; // @[Cat.scala 31:58]
  wire [15:0] canValid_lo = {_canValid_T_33,_canValid_T_35,_canValid_T_37,_canValid_T_39,_canValid_T_41,_canValid_T_43,
    _canValid_T_45,_canValid_T_47,canValid_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] canValid_hi_lo = {_canValid_T_17,_canValid_T_19,_canValid_T_21,_canValid_T_23,_canValid_T_25,_canValid_T_27
    ,_canValid_T_29,_canValid_T_31}; // @[Cat.scala 31:58]
  wire [31:0] _canValid_T_64 = {_canValid_T_1,_canValid_T_3,_canValid_T_5,_canValid_T_7,_canValid_T_9,_canValid_T_11,
    _canValid_T_13,_canValid_T_15,canValid_hi_lo,canValid_lo}; // @[Cat.scala 31:58]
  wire  _T_400 = io_validResp_out_ready & io_validResp_out_valid; // @[Decoupled.scala 50:35]
  wire [4:0] rspIdx = io_validResp_out_bits_source[18:14]; // @[WriteStack.scala 166:48]
  wire [1:0] _GEN_1280 = 5'h0 == rspIdx ? 2'h3 : _GEN_1216; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1281 = 5'h1 == rspIdx ? 2'h3 : _GEN_1218; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1282 = 5'h2 == rspIdx ? 2'h3 : _GEN_1220; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1283 = 5'h3 == rspIdx ? 2'h3 : _GEN_1222; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1284 = 5'h4 == rspIdx ? 2'h3 : _GEN_1224; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1285 = 5'h5 == rspIdx ? 2'h3 : _GEN_1226; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1286 = 5'h6 == rspIdx ? 2'h3 : _GEN_1228; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1287 = 5'h7 == rspIdx ? 2'h3 : _GEN_1230; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1288 = 5'h8 == rspIdx ? 2'h3 : _GEN_1232; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1289 = 5'h9 == rspIdx ? 2'h3 : _GEN_1234; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1290 = 5'ha == rspIdx ? 2'h3 : _GEN_1236; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1291 = 5'hb == rspIdx ? 2'h3 : _GEN_1238; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1292 = 5'hc == rspIdx ? 2'h3 : _GEN_1240; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1293 = 5'hd == rspIdx ? 2'h3 : _GEN_1242; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1294 = 5'he == rspIdx ? 2'h3 : _GEN_1244; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1295 = 5'hf == rspIdx ? 2'h3 : _GEN_1246; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1296 = 5'h10 == rspIdx ? 2'h3 : _GEN_1248; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1297 = 5'h11 == rspIdx ? 2'h3 : _GEN_1250; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1298 = 5'h12 == rspIdx ? 2'h3 : _GEN_1252; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1299 = 5'h13 == rspIdx ? 2'h3 : _GEN_1254; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1300 = 5'h14 == rspIdx ? 2'h3 : _GEN_1256; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1301 = 5'h15 == rspIdx ? 2'h3 : _GEN_1258; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1302 = 5'h16 == rspIdx ? 2'h3 : _GEN_1260; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1303 = 5'h17 == rspIdx ? 2'h3 : _GEN_1262; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1304 = 5'h18 == rspIdx ? 2'h3 : _GEN_1264; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1305 = 5'h19 == rspIdx ? 2'h3 : _GEN_1266; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1306 = 5'h1a == rspIdx ? 2'h3 : _GEN_1268; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1307 = 5'h1b == rspIdx ? 2'h3 : _GEN_1270; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1308 = 5'h1c == rspIdx ? 2'h3 : _GEN_1272; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1309 = 5'h1d == rspIdx ? 2'h3 : _GEN_1274; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1310 = 5'h1e == rspIdx ? 2'h3 : _GEN_1276; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1311 = 5'h1f == rspIdx ? 2'h3 : _GEN_1278; // @[WriteStack.scala 168:{25,25}]
  wire [1:0] _GEN_1312 = _T_400 ? _GEN_1280 : _GEN_1216; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1313 = _T_400 ? _GEN_1281 : _GEN_1218; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1314 = _T_400 ? _GEN_1282 : _GEN_1220; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1315 = _T_400 ? _GEN_1283 : _GEN_1222; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1316 = _T_400 ? _GEN_1284 : _GEN_1224; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1317 = _T_400 ? _GEN_1285 : _GEN_1226; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1318 = _T_400 ? _GEN_1286 : _GEN_1228; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1319 = _T_400 ? _GEN_1287 : _GEN_1230; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1320 = _T_400 ? _GEN_1288 : _GEN_1232; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1321 = _T_400 ? _GEN_1289 : _GEN_1234; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1322 = _T_400 ? _GEN_1290 : _GEN_1236; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1323 = _T_400 ? _GEN_1291 : _GEN_1238; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1324 = _T_400 ? _GEN_1292 : _GEN_1240; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1325 = _T_400 ? _GEN_1293 : _GEN_1242; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1326 = _T_400 ? _GEN_1294 : _GEN_1244; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1327 = _T_400 ? _GEN_1295 : _GEN_1246; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1328 = _T_400 ? _GEN_1296 : _GEN_1248; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1329 = _T_400 ? _GEN_1297 : _GEN_1250; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1330 = _T_400 ? _GEN_1298 : _GEN_1252; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1331 = _T_400 ? _GEN_1299 : _GEN_1254; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1332 = _T_400 ? _GEN_1300 : _GEN_1256; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1333 = _T_400 ? _GEN_1301 : _GEN_1258; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1334 = _T_400 ? _GEN_1302 : _GEN_1260; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1335 = _T_400 ? _GEN_1303 : _GEN_1262; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1336 = _T_400 ? _GEN_1304 : _GEN_1264; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1337 = _T_400 ? _GEN_1305 : _GEN_1266; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1338 = _T_400 ? _GEN_1306 : _GEN_1268; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1339 = _T_400 ? _GEN_1307 : _GEN_1270; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1340 = _T_400 ? _GEN_1308 : _GEN_1272; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1341 = _T_400 ? _GEN_1309 : _GEN_1274; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1342 = _T_400 ? _GEN_1310 : _GEN_1276; // @[WriteStack.scala 165:5]
  wire [1:0] _GEN_1343 = _T_400 ? _GEN_1311 : _GEN_1278; // @[WriteStack.scala 165:5]
  wire  _canAW_T = _GEN_1856 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_2 = writeStack_0_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_3 = writeStack_0_wvalid & _GEN_1856 == 3'h2 & writeStack_0_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_4 = writeStack_0_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_5 = writeStack_0_wvalid & _GEN_1856 == 3'h2 & writeStack_0_validStatus == 2'h3 &
    writeStack_0_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_6 = _GEN_1857 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_8 = writeStack_1_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_9 = writeStack_1_wvalid & _GEN_1857 == 3'h2 & writeStack_1_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_10 = writeStack_1_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_11 = writeStack_1_wvalid & _GEN_1857 == 3'h2 & writeStack_1_validStatus == 2'h3 &
    writeStack_1_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_12 = _GEN_1858 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_14 = writeStack_2_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_15 = writeStack_2_wvalid & _GEN_1858 == 3'h2 & writeStack_2_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_16 = writeStack_2_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_17 = writeStack_2_wvalid & _GEN_1858 == 3'h2 & writeStack_2_validStatus == 2'h3 &
    writeStack_2_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_18 = _GEN_1859 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_20 = writeStack_3_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_21 = writeStack_3_wvalid & _GEN_1859 == 3'h2 & writeStack_3_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_22 = writeStack_3_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_23 = writeStack_3_wvalid & _GEN_1859 == 3'h2 & writeStack_3_validStatus == 2'h3 &
    writeStack_3_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_24 = _GEN_1860 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_26 = writeStack_4_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_27 = writeStack_4_wvalid & _GEN_1860 == 3'h2 & writeStack_4_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_28 = writeStack_4_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_29 = writeStack_4_wvalid & _GEN_1860 == 3'h2 & writeStack_4_validStatus == 2'h3 &
    writeStack_4_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_30 = _GEN_1861 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_32 = writeStack_5_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_33 = writeStack_5_wvalid & _GEN_1861 == 3'h2 & writeStack_5_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_34 = writeStack_5_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_35 = writeStack_5_wvalid & _GEN_1861 == 3'h2 & writeStack_5_validStatus == 2'h3 &
    writeStack_5_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_36 = _GEN_1862 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_38 = writeStack_6_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_39 = writeStack_6_wvalid & _GEN_1862 == 3'h2 & writeStack_6_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_40 = writeStack_6_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_41 = writeStack_6_wvalid & _GEN_1862 == 3'h2 & writeStack_6_validStatus == 2'h3 &
    writeStack_6_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_42 = _GEN_1863 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_44 = writeStack_7_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_45 = writeStack_7_wvalid & _GEN_1863 == 3'h2 & writeStack_7_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_46 = writeStack_7_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_47 = writeStack_7_wvalid & _GEN_1863 == 3'h2 & writeStack_7_validStatus == 2'h3 &
    writeStack_7_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_48 = _GEN_1864 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_50 = writeStack_8_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_51 = writeStack_8_wvalid & _GEN_1864 == 3'h2 & writeStack_8_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_52 = writeStack_8_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_53 = writeStack_8_wvalid & _GEN_1864 == 3'h2 & writeStack_8_validStatus == 2'h3 &
    writeStack_8_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_54 = _GEN_1865 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_56 = writeStack_9_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_57 = writeStack_9_wvalid & _GEN_1865 == 3'h2 & writeStack_9_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_58 = writeStack_9_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_59 = writeStack_9_wvalid & _GEN_1865 == 3'h2 & writeStack_9_validStatus == 2'h3 &
    writeStack_9_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_60 = _GEN_1866 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_62 = writeStack_10_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_63 = writeStack_10_wvalid & _GEN_1866 == 3'h2 & writeStack_10_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_64 = writeStack_10_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_65 = writeStack_10_wvalid & _GEN_1866 == 3'h2 & writeStack_10_validStatus == 2'h3 &
    writeStack_10_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_66 = _GEN_1867 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_68 = writeStack_11_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_69 = writeStack_11_wvalid & _GEN_1867 == 3'h2 & writeStack_11_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_70 = writeStack_11_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_71 = writeStack_11_wvalid & _GEN_1867 == 3'h2 & writeStack_11_validStatus == 2'h3 &
    writeStack_11_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_72 = _GEN_1868 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_74 = writeStack_12_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_75 = writeStack_12_wvalid & _GEN_1868 == 3'h2 & writeStack_12_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_76 = writeStack_12_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_77 = writeStack_12_wvalid & _GEN_1868 == 3'h2 & writeStack_12_validStatus == 2'h3 &
    writeStack_12_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_78 = _GEN_1869 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_80 = writeStack_13_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_81 = writeStack_13_wvalid & _GEN_1869 == 3'h2 & writeStack_13_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_82 = writeStack_13_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_83 = writeStack_13_wvalid & _GEN_1869 == 3'h2 & writeStack_13_validStatus == 2'h3 &
    writeStack_13_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_84 = _GEN_1870 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_86 = writeStack_14_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_87 = writeStack_14_wvalid & _GEN_1870 == 3'h2 & writeStack_14_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_88 = writeStack_14_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_89 = writeStack_14_wvalid & _GEN_1870 == 3'h2 & writeStack_14_validStatus == 2'h3 &
    writeStack_14_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_90 = _GEN_1871 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_92 = writeStack_15_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_93 = writeStack_15_wvalid & _GEN_1871 == 3'h2 & writeStack_15_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_94 = writeStack_15_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_95 = writeStack_15_wvalid & _GEN_1871 == 3'h2 & writeStack_15_validStatus == 2'h3 &
    writeStack_15_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_96 = _GEN_1872 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_98 = writeStack_16_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_99 = writeStack_16_wvalid & _GEN_1872 == 3'h2 & writeStack_16_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_100 = writeStack_16_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_101 = writeStack_16_wvalid & _GEN_1872 == 3'h2 & writeStack_16_validStatus == 2'h3 &
    writeStack_16_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_102 = _GEN_1873 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_104 = writeStack_17_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_105 = writeStack_17_wvalid & _GEN_1873 == 3'h2 & writeStack_17_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_106 = writeStack_17_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_107 = writeStack_17_wvalid & _GEN_1873 == 3'h2 & writeStack_17_validStatus == 2'h3 &
    writeStack_17_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_108 = _GEN_1874 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_110 = writeStack_18_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_111 = writeStack_18_wvalid & _GEN_1874 == 3'h2 & writeStack_18_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_112 = writeStack_18_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_113 = writeStack_18_wvalid & _GEN_1874 == 3'h2 & writeStack_18_validStatus == 2'h3 &
    writeStack_18_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_114 = _GEN_1875 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_116 = writeStack_19_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_117 = writeStack_19_wvalid & _GEN_1875 == 3'h2 & writeStack_19_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_118 = writeStack_19_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_119 = writeStack_19_wvalid & _GEN_1875 == 3'h2 & writeStack_19_validStatus == 2'h3 &
    writeStack_19_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_120 = _GEN_1876 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_122 = writeStack_20_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_123 = writeStack_20_wvalid & _GEN_1876 == 3'h2 & writeStack_20_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_124 = writeStack_20_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_125 = writeStack_20_wvalid & _GEN_1876 == 3'h2 & writeStack_20_validStatus == 2'h3 &
    writeStack_20_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_126 = _GEN_1877 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_128 = writeStack_21_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_129 = writeStack_21_wvalid & _GEN_1877 == 3'h2 & writeStack_21_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_130 = writeStack_21_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_131 = writeStack_21_wvalid & _GEN_1877 == 3'h2 & writeStack_21_validStatus == 2'h3 &
    writeStack_21_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_132 = _GEN_1878 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_134 = writeStack_22_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_135 = writeStack_22_wvalid & _GEN_1878 == 3'h2 & writeStack_22_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_136 = writeStack_22_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_137 = writeStack_22_wvalid & _GEN_1878 == 3'h2 & writeStack_22_validStatus == 2'h3 &
    writeStack_22_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_138 = _GEN_1879 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_140 = writeStack_23_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_141 = writeStack_23_wvalid & _GEN_1879 == 3'h2 & writeStack_23_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_142 = writeStack_23_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_143 = writeStack_23_wvalid & _GEN_1879 == 3'h2 & writeStack_23_validStatus == 2'h3 &
    writeStack_23_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_144 = _GEN_1880 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_146 = writeStack_24_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_147 = writeStack_24_wvalid & _GEN_1880 == 3'h2 & writeStack_24_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_148 = writeStack_24_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_149 = writeStack_24_wvalid & _GEN_1880 == 3'h2 & writeStack_24_validStatus == 2'h3 &
    writeStack_24_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_150 = _GEN_1881 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_152 = writeStack_25_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_153 = writeStack_25_wvalid & _GEN_1881 == 3'h2 & writeStack_25_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_154 = writeStack_25_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_155 = writeStack_25_wvalid & _GEN_1881 == 3'h2 & writeStack_25_validStatus == 2'h3 &
    writeStack_25_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_156 = _GEN_1882 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_158 = writeStack_26_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_159 = writeStack_26_wvalid & _GEN_1882 == 3'h2 & writeStack_26_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_160 = writeStack_26_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_161 = writeStack_26_wvalid & _GEN_1882 == 3'h2 & writeStack_26_validStatus == 2'h3 &
    writeStack_26_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_162 = _GEN_1883 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_164 = writeStack_27_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_165 = writeStack_27_wvalid & _GEN_1883 == 3'h2 & writeStack_27_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_166 = writeStack_27_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_167 = writeStack_27_wvalid & _GEN_1883 == 3'h2 & writeStack_27_validStatus == 2'h3 &
    writeStack_27_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_168 = _GEN_1884 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_170 = writeStack_28_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_171 = writeStack_28_wvalid & _GEN_1884 == 3'h2 & writeStack_28_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_172 = writeStack_28_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_173 = writeStack_28_wvalid & _GEN_1884 == 3'h2 & writeStack_28_validStatus == 2'h3 &
    writeStack_28_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_174 = _GEN_1885 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_176 = writeStack_29_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_177 = writeStack_29_wvalid & _GEN_1885 == 3'h2 & writeStack_29_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_178 = writeStack_29_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_179 = writeStack_29_wvalid & _GEN_1885 == 3'h2 & writeStack_29_validStatus == 2'h3 &
    writeStack_29_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_180 = _GEN_1886 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_182 = writeStack_30_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_183 = writeStack_30_wvalid & _GEN_1886 == 3'h2 & writeStack_30_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_184 = writeStack_30_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_185 = writeStack_30_wvalid & _GEN_1886 == 3'h2 & writeStack_30_validStatus == 2'h3 &
    writeStack_30_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _canAW_T_186 = _GEN_1887 == 3'h2; // @[WriteStack.scala 173:61]
  wire  _canAW_T_188 = writeStack_31_validStatus == 2'h3; // @[WriteStack.scala 173:89]
  wire  _canAW_T_189 = writeStack_31_wvalid & _GEN_1887 == 3'h2 & writeStack_31_validStatus == 2'h3; // @[WriteStack.scala 173:73]
  wire  _canAW_T_190 = writeStack_31_entryFifoid == 5'h0; // @[WriteStack.scala 173:120]
  wire  _canAW_T_191 = writeStack_31_wvalid & _GEN_1887 == 3'h2 & writeStack_31_validStatus == 2'h3 &
    writeStack_31_entryFifoid == 5'h0; // @[WriteStack.scala 173:103]
  wire  _T_402 = io_axiMenWriteReq_out_w_ready & io_axiMenWriteReq_out_w_valid; // @[Decoupled.scala 50:35]
  wire  _T_403 = _T & _T_402; // @[WriteStack.scala 193:34]
  wire  _writeStack_entryFifoid_T_3 = _GEN_1856 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_5 = writeStack_0_wvalid & (_canW_T | _canAW_T | _GEN_1856 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_9 = _GEN_1857 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_11 = writeStack_1_wvalid & (_canW_T_4 | _canAW_T_6 | _GEN_1857 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_15 = _GEN_1858 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_17 = writeStack_2_wvalid & (_canW_T_8 | _canAW_T_12 | _GEN_1858 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_21 = _GEN_1859 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_23 = writeStack_3_wvalid & (_canW_T_12 | _canAW_T_18 | _GEN_1859 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_27 = _GEN_1860 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_29 = writeStack_4_wvalid & (_canW_T_16 | _canAW_T_24 | _GEN_1860 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_33 = _GEN_1861 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_35 = writeStack_5_wvalid & (_canW_T_20 | _canAW_T_30 | _GEN_1861 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_39 = _GEN_1862 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_41 = writeStack_6_wvalid & (_canW_T_24 | _canAW_T_36 | _GEN_1862 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_45 = _GEN_1863 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_47 = writeStack_7_wvalid & (_canW_T_28 | _canAW_T_42 | _GEN_1863 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_51 = _GEN_1864 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_53 = writeStack_8_wvalid & (_canW_T_32 | _canAW_T_48 | _GEN_1864 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_57 = _GEN_1865 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_59 = writeStack_9_wvalid & (_canW_T_36 | _canAW_T_54 | _GEN_1865 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_63 = _GEN_1866 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_65 = writeStack_10_wvalid & (_canW_T_40 | _canAW_T_60 | _GEN_1866 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_69 = _GEN_1867 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_71 = writeStack_11_wvalid & (_canW_T_44 | _canAW_T_66 | _GEN_1867 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_75 = _GEN_1868 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_77 = writeStack_12_wvalid & (_canW_T_48 | _canAW_T_72 | _GEN_1868 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_81 = _GEN_1869 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_83 = writeStack_13_wvalid & (_canW_T_52 | _canAW_T_78 | _GEN_1869 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_87 = _GEN_1870 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_89 = writeStack_14_wvalid & (_canW_T_56 | _canAW_T_84 | _GEN_1870 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_93 = _GEN_1871 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_95 = writeStack_15_wvalid & (_canW_T_60 | _canAW_T_90 | _GEN_1871 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_99 = _GEN_1872 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_101 = writeStack_16_wvalid & (_canW_T_64 | _canAW_T_96 | _GEN_1872 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_105 = _GEN_1873 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_107 = writeStack_17_wvalid & (_canW_T_68 | _canAW_T_102 | _GEN_1873 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_111 = _GEN_1874 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_113 = writeStack_18_wvalid & (_canW_T_72 | _canAW_T_108 | _GEN_1874 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_117 = _GEN_1875 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_119 = writeStack_19_wvalid & (_canW_T_76 | _canAW_T_114 | _GEN_1875 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_123 = _GEN_1876 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_125 = writeStack_20_wvalid & (_canW_T_80 | _canAW_T_120 | _GEN_1876 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_129 = _GEN_1877 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_131 = writeStack_21_wvalid & (_canW_T_84 | _canAW_T_126 | _GEN_1877 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_135 = _GEN_1878 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_137 = writeStack_22_wvalid & (_canW_T_88 | _canAW_T_132 | _GEN_1878 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_141 = _GEN_1879 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_143 = writeStack_23_wvalid & (_canW_T_92 | _canAW_T_138 | _GEN_1879 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_147 = _GEN_1880 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_149 = writeStack_24_wvalid & (_canW_T_96 | _canAW_T_144 | _GEN_1880 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_153 = _GEN_1881 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_155 = writeStack_25_wvalid & (_canW_T_100 | _canAW_T_150 | _GEN_1881 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_159 = _GEN_1882 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_161 = writeStack_26_wvalid & (_canW_T_104 | _canAW_T_156 | _GEN_1882 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_165 = _GEN_1883 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_167 = writeStack_27_wvalid & (_canW_T_108 | _canAW_T_162 | _GEN_1883 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_171 = _GEN_1884 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_173 = writeStack_28_wvalid & (_canW_T_112 | _canAW_T_168 | _GEN_1884 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_177 = _GEN_1885 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_179 = writeStack_29_wvalid & (_canW_T_116 | _canAW_T_174 | _GEN_1885 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_183 = _GEN_1886 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_185 = writeStack_30_wvalid & (_canW_T_120 | _canAW_T_180 | _GEN_1886 == 3'h3); // @[WriteStack.scala 196:64]
  wire  _writeStack_entryFifoid_T_189 = _GEN_1887 == 3'h3; // @[WriteStack.scala 196:126]
  wire  _writeStack_entryFifoid_T_191 = writeStack_31_wvalid & (_canW_T_124 | _canAW_T_186 | _GEN_1887 == 3'h3); // @[WriteStack.scala 196:64]
  wire [1:0] _writeStack_entryFifoid_T_192 = _writeStack_entryFifoid_T_5 + _writeStack_entryFifoid_T_11; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_194 = _writeStack_entryFifoid_T_17 + _writeStack_entryFifoid_T_23; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_196 = _writeStack_entryFifoid_T_192 + _writeStack_entryFifoid_T_194; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_198 = _writeStack_entryFifoid_T_29 + _writeStack_entryFifoid_T_35; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_200 = _writeStack_entryFifoid_T_41 + _writeStack_entryFifoid_T_47; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_202 = _writeStack_entryFifoid_T_198 + _writeStack_entryFifoid_T_200; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_entryFifoid_T_204 = _writeStack_entryFifoid_T_196 + _writeStack_entryFifoid_T_202; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_206 = _writeStack_entryFifoid_T_53 + _writeStack_entryFifoid_T_59; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_208 = _writeStack_entryFifoid_T_65 + _writeStack_entryFifoid_T_71; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_210 = _writeStack_entryFifoid_T_206 + _writeStack_entryFifoid_T_208; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_212 = _writeStack_entryFifoid_T_77 + _writeStack_entryFifoid_T_83; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_214 = _writeStack_entryFifoid_T_89 + _writeStack_entryFifoid_T_95; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_216 = _writeStack_entryFifoid_T_212 + _writeStack_entryFifoid_T_214; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_entryFifoid_T_218 = _writeStack_entryFifoid_T_210 + _writeStack_entryFifoid_T_216; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_entryFifoid_T_220 = _writeStack_entryFifoid_T_204 + _writeStack_entryFifoid_T_218; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_222 = _writeStack_entryFifoid_T_101 + _writeStack_entryFifoid_T_107; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_224 = _writeStack_entryFifoid_T_113 + _writeStack_entryFifoid_T_119; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_226 = _writeStack_entryFifoid_T_222 + _writeStack_entryFifoid_T_224; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_228 = _writeStack_entryFifoid_T_125 + _writeStack_entryFifoid_T_131; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_230 = _writeStack_entryFifoid_T_137 + _writeStack_entryFifoid_T_143; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_232 = _writeStack_entryFifoid_T_228 + _writeStack_entryFifoid_T_230; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_entryFifoid_T_234 = _writeStack_entryFifoid_T_226 + _writeStack_entryFifoid_T_232; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_236 = _writeStack_entryFifoid_T_149 + _writeStack_entryFifoid_T_155; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_238 = _writeStack_entryFifoid_T_161 + _writeStack_entryFifoid_T_167; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_240 = _writeStack_entryFifoid_T_236 + _writeStack_entryFifoid_T_238; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_242 = _writeStack_entryFifoid_T_173 + _writeStack_entryFifoid_T_179; // @[Bitwise.scala 48:55]
  wire [1:0] _writeStack_entryFifoid_T_244 = _writeStack_entryFifoid_T_185 + _writeStack_entryFifoid_T_191; // @[Bitwise.scala 48:55]
  wire [2:0] _writeStack_entryFifoid_T_246 = _writeStack_entryFifoid_T_242 + _writeStack_entryFifoid_T_244; // @[Bitwise.scala 48:55]
  wire [3:0] _writeStack_entryFifoid_T_248 = _writeStack_entryFifoid_T_240 + _writeStack_entryFifoid_T_246; // @[Bitwise.scala 48:55]
  wire [4:0] _writeStack_entryFifoid_T_250 = _writeStack_entryFifoid_T_234 + _writeStack_entryFifoid_T_248; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_entryFifoid_T_252 = _writeStack_entryFifoid_T_220 + _writeStack_entryFifoid_T_250; // @[Bitwise.scala 48:55]
  wire [5:0] _writeStack_entryFifoid_T_255 = _writeStack_entryFifoid_T_252 - 6'h1; // @[WriteStack.scala 196:139]
  wire [4:0] _GEN_1344 = 5'h0 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_0_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1345 = 5'h1 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_1_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1346 = 5'h2 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_2_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1347 = 5'h3 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_3_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1348 = 5'h4 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_4_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1349 = 5'h5 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_5_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1350 = 5'h6 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_6_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1351 = 5'h7 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_7_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1352 = 5'h8 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_8_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1353 = 5'h9 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_9_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1354 = 5'ha == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_10_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1355 = 5'hb == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_11_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1356 = 5'hc == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_12_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1357 = 5'hd == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_13_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1358 = 5'he == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_14_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1359 = 5'hf == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_15_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1360 = 5'h10 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_16_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1361 = 5'h11 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_17_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1362 = 5'h12 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_18_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1363 = 5'h13 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_19_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1364 = 5'h14 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_20_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1365 = 5'h15 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_21_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1366 = 5'h16 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_22_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1367 = 5'h17 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_23_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1368 = 5'h18 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_24_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1369 = 5'h19 == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_25_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1370 = 5'h1a == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_26_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1371 = 5'h1b == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_27_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1372 = 5'h1c == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_28_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1373 = 5'h1d == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_29_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1374 = 5'h1e == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_30_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire [4:0] _GEN_1375 = 5'h1f == idxInsert ? _writeStack_entryFifoid_T_255[4:0] : writeStack_31_entryFifoid; // @[WriteStack.scala 196:{23,23} 56:27]
  wire  _T_407 = _T & ~_T_402; // @[WriteStack.scala 197:40]
  wire [4:0] _GEN_1376 = 5'h0 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_0_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1377 = 5'h1 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_1_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1378 = 5'h2 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_2_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1379 = 5'h3 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_3_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1380 = 5'h4 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_4_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1381 = 5'h5 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_5_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1382 = 5'h6 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_6_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1383 = 5'h7 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_7_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1384 = 5'h8 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_8_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1385 = 5'h9 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_9_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1386 = 5'ha == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_10_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1387 = 5'hb == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_11_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1388 = 5'hc == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_12_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1389 = 5'hd == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_13_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1390 = 5'he == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_14_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1391 = 5'hf == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_15_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1392 = 5'h10 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_16_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1393 = 5'h11 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_17_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1394 = 5'h12 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_18_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1395 = 5'h13 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_19_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1396 = 5'h14 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_20_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1397 = 5'h15 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_21_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1398 = 5'h16 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_22_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1399 = 5'h17 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_23_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1400 = 5'h18 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_24_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1401 = 5'h19 == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_25_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1402 = 5'h1a == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_26_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1403 = 5'h1b == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_27_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1404 = 5'h1c == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_28_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1405 = 5'h1d == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_29_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1406 = 5'h1e == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_30_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1407 = 5'h1f == idxInsert ? _writeStack_entryFifoid_T_252[4:0] : writeStack_31_entryFifoid; // @[WriteStack.scala 200:{23,23} 56:27]
  wire [4:0] _GEN_1408 = _T_407 ? _GEN_1376 : writeStack_0_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1409 = _T_407 ? _GEN_1377 : writeStack_1_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1410 = _T_407 ? _GEN_1378 : writeStack_2_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1411 = _T_407 ? _GEN_1379 : writeStack_3_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1412 = _T_407 ? _GEN_1380 : writeStack_4_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1413 = _T_407 ? _GEN_1381 : writeStack_5_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1414 = _T_407 ? _GEN_1382 : writeStack_6_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1415 = _T_407 ? _GEN_1383 : writeStack_7_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1416 = _T_407 ? _GEN_1384 : writeStack_8_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1417 = _T_407 ? _GEN_1385 : writeStack_9_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1418 = _T_407 ? _GEN_1386 : writeStack_10_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1419 = _T_407 ? _GEN_1387 : writeStack_11_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1420 = _T_407 ? _GEN_1388 : writeStack_12_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1421 = _T_407 ? _GEN_1389 : writeStack_13_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1422 = _T_407 ? _GEN_1390 : writeStack_14_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1423 = _T_407 ? _GEN_1391 : writeStack_15_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1424 = _T_407 ? _GEN_1392 : writeStack_16_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1425 = _T_407 ? _GEN_1393 : writeStack_17_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1426 = _T_407 ? _GEN_1394 : writeStack_18_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1427 = _T_407 ? _GEN_1395 : writeStack_19_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1428 = _T_407 ? _GEN_1396 : writeStack_20_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1429 = _T_407 ? _GEN_1397 : writeStack_21_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1430 = _T_407 ? _GEN_1398 : writeStack_22_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1431 = _T_407 ? _GEN_1399 : writeStack_23_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1432 = _T_407 ? _GEN_1400 : writeStack_24_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1433 = _T_407 ? _GEN_1401 : writeStack_25_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1434 = _T_407 ? _GEN_1402 : writeStack_26_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1435 = _T_407 ? _GEN_1403 : writeStack_27_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1436 = _T_407 ? _GEN_1404 : writeStack_28_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1437 = _T_407 ? _GEN_1405 : writeStack_29_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1438 = _T_407 ? _GEN_1406 : writeStack_30_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1439 = _T_407 ? _GEN_1407 : writeStack_31_entryFifoid; // @[WriteStack.scala 198:3 56:27]
  wire [4:0] _GEN_1440 = _T_403 ? _GEN_1344 : _GEN_1408; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1441 = _T_403 ? _GEN_1345 : _GEN_1409; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1442 = _T_403 ? _GEN_1346 : _GEN_1410; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1443 = _T_403 ? _GEN_1347 : _GEN_1411; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1444 = _T_403 ? _GEN_1348 : _GEN_1412; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1445 = _T_403 ? _GEN_1349 : _GEN_1413; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1446 = _T_403 ? _GEN_1350 : _GEN_1414; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1447 = _T_403 ? _GEN_1351 : _GEN_1415; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1448 = _T_403 ? _GEN_1352 : _GEN_1416; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1449 = _T_403 ? _GEN_1353 : _GEN_1417; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1450 = _T_403 ? _GEN_1354 : _GEN_1418; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1451 = _T_403 ? _GEN_1355 : _GEN_1419; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1452 = _T_403 ? _GEN_1356 : _GEN_1420; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1453 = _T_403 ? _GEN_1357 : _GEN_1421; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1454 = _T_403 ? _GEN_1358 : _GEN_1422; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1455 = _T_403 ? _GEN_1359 : _GEN_1423; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1456 = _T_403 ? _GEN_1360 : _GEN_1424; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1457 = _T_403 ? _GEN_1361 : _GEN_1425; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1458 = _T_403 ? _GEN_1362 : _GEN_1426; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1459 = _T_403 ? _GEN_1363 : _GEN_1427; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1460 = _T_403 ? _GEN_1364 : _GEN_1428; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1461 = _T_403 ? _GEN_1365 : _GEN_1429; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1462 = _T_403 ? _GEN_1366 : _GEN_1430; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1463 = _T_403 ? _GEN_1367 : _GEN_1431; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1464 = _T_403 ? _GEN_1368 : _GEN_1432; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1465 = _T_403 ? _GEN_1369 : _GEN_1433; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1466 = _T_403 ? _GEN_1370 : _GEN_1434; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1467 = _T_403 ? _GEN_1371 : _GEN_1435; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1468 = _T_403 ? _GEN_1372 : _GEN_1436; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1469 = _T_403 ? _GEN_1373 : _GEN_1437; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1470 = _T_403 ? _GEN_1374 : _GEN_1438; // @[WriteStack.scala 194:3]
  wire [4:0] _GEN_1471 = _T_403 ? _GEN_1375 : _GEN_1439; // @[WriteStack.scala 194:3]
  wire  _T_408 = io_axiMenWriteReq_out_aw_ready & io_axiMenWriteReq_out_aw_valid; // @[Decoupled.scala 50:35]
  wire [2:0] _GEN_1472 = _canAW_T_5 ? 3'h3 : _GEN_866; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1473 = _canAW_T_11 ? 3'h3 : _GEN_870; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1474 = _canAW_T_17 ? 3'h3 : _GEN_874; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1475 = _canAW_T_23 ? 3'h3 : _GEN_878; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1476 = _canAW_T_29 ? 3'h3 : _GEN_882; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1477 = _canAW_T_35 ? 3'h3 : _GEN_886; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1478 = _canAW_T_41 ? 3'h3 : _GEN_890; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1479 = _canAW_T_47 ? 3'h3 : _GEN_894; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1480 = _canAW_T_53 ? 3'h3 : _GEN_898; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1481 = _canAW_T_59 ? 3'h3 : _GEN_902; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1482 = _canAW_T_65 ? 3'h3 : _GEN_906; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1483 = _canAW_T_71 ? 3'h3 : _GEN_910; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1484 = _canAW_T_77 ? 3'h3 : _GEN_914; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1485 = _canAW_T_83 ? 3'h3 : _GEN_918; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1486 = _canAW_T_89 ? 3'h3 : _GEN_922; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1487 = _canAW_T_95 ? 3'h3 : _GEN_926; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1488 = _canAW_T_101 ? 3'h3 : _GEN_930; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1489 = _canAW_T_107 ? 3'h3 : _GEN_934; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1490 = _canAW_T_113 ? 3'h3 : _GEN_938; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1491 = _canAW_T_119 ? 3'h3 : _GEN_942; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1492 = _canAW_T_125 ? 3'h3 : _GEN_946; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1493 = _canAW_T_131 ? 3'h3 : _GEN_950; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1494 = _canAW_T_137 ? 3'h3 : _GEN_954; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1495 = _canAW_T_143 ? 3'h3 : _GEN_958; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1496 = _canAW_T_149 ? 3'h3 : _GEN_962; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1497 = _canAW_T_155 ? 3'h3 : _GEN_966; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1498 = _canAW_T_161 ? 3'h3 : _GEN_970; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1499 = _canAW_T_167 ? 3'h3 : _GEN_974; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1500 = _canAW_T_173 ? 3'h3 : _GEN_978; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1501 = _canAW_T_179 ? 3'h3 : _GEN_982; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1502 = _canAW_T_185 ? 3'h3 : _GEN_986; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1503 = _canAW_T_191 ? 3'h3 : _GEN_990; // @[WriteStack.scala 207:17 209:31]
  wire [2:0] _GEN_1504 = _T_408 ? _GEN_1472 : _GEN_866; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1505 = _T_408 ? _GEN_1473 : _GEN_870; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1506 = _T_408 ? _GEN_1474 : _GEN_874; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1507 = _T_408 ? _GEN_1475 : _GEN_878; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1508 = _T_408 ? _GEN_1476 : _GEN_882; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1509 = _T_408 ? _GEN_1477 : _GEN_886; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1510 = _T_408 ? _GEN_1478 : _GEN_890; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1511 = _T_408 ? _GEN_1479 : _GEN_894; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1512 = _T_408 ? _GEN_1480 : _GEN_898; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1513 = _T_408 ? _GEN_1481 : _GEN_902; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1514 = _T_408 ? _GEN_1482 : _GEN_906; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1515 = _T_408 ? _GEN_1483 : _GEN_910; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1516 = _T_408 ? _GEN_1484 : _GEN_914; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1517 = _T_408 ? _GEN_1485 : _GEN_918; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1518 = _T_408 ? _GEN_1486 : _GEN_922; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1519 = _T_408 ? _GEN_1487 : _GEN_926; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1520 = _T_408 ? _GEN_1488 : _GEN_930; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1521 = _T_408 ? _GEN_1489 : _GEN_934; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1522 = _T_408 ? _GEN_1490 : _GEN_938; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1523 = _T_408 ? _GEN_1491 : _GEN_942; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1524 = _T_408 ? _GEN_1492 : _GEN_946; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1525 = _T_408 ? _GEN_1493 : _GEN_950; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1526 = _T_408 ? _GEN_1494 : _GEN_954; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1527 = _T_408 ? _GEN_1495 : _GEN_958; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1528 = _T_408 ? _GEN_1496 : _GEN_962; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1529 = _T_408 ? _GEN_1497 : _GEN_966; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1530 = _T_408 ? _GEN_1498 : _GEN_970; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1531 = _T_408 ? _GEN_1499 : _GEN_974; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1532 = _T_408 ? _GEN_1500 : _GEN_978; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1533 = _T_408 ? _GEN_1501 : _GEN_982; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1534 = _T_408 ? _GEN_1502 : _GEN_986; // @[WriteStack.scala 203:5]
  wire [2:0] _GEN_1535 = _T_408 ? _GEN_1503 : _GEN_990; // @[WriteStack.scala 203:5]
  wire  _canMenW_T_3 = writeStack_0_wvalid & _writeStack_entryFifoid_T_3 & _canAW_T_2; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_5 = writeStack_0_wvalid & _writeStack_entryFifoid_T_3 & _canAW_T_2 & _canAW_T_4; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_9 = writeStack_1_wvalid & _writeStack_entryFifoid_T_9 & _canAW_T_8; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_11 = writeStack_1_wvalid & _writeStack_entryFifoid_T_9 & _canAW_T_8 & _canAW_T_10; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_15 = writeStack_2_wvalid & _writeStack_entryFifoid_T_15 & _canAW_T_14; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_17 = writeStack_2_wvalid & _writeStack_entryFifoid_T_15 & _canAW_T_14 & _canAW_T_16; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_21 = writeStack_3_wvalid & _writeStack_entryFifoid_T_21 & _canAW_T_20; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_23 = writeStack_3_wvalid & _writeStack_entryFifoid_T_21 & _canAW_T_20 & _canAW_T_22; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_27 = writeStack_4_wvalid & _writeStack_entryFifoid_T_27 & _canAW_T_26; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_29 = writeStack_4_wvalid & _writeStack_entryFifoid_T_27 & _canAW_T_26 & _canAW_T_28; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_33 = writeStack_5_wvalid & _writeStack_entryFifoid_T_33 & _canAW_T_32; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_35 = writeStack_5_wvalid & _writeStack_entryFifoid_T_33 & _canAW_T_32 & _canAW_T_34; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_39 = writeStack_6_wvalid & _writeStack_entryFifoid_T_39 & _canAW_T_38; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_41 = writeStack_6_wvalid & _writeStack_entryFifoid_T_39 & _canAW_T_38 & _canAW_T_40; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_45 = writeStack_7_wvalid & _writeStack_entryFifoid_T_45 & _canAW_T_44; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_47 = writeStack_7_wvalid & _writeStack_entryFifoid_T_45 & _canAW_T_44 & _canAW_T_46; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_51 = writeStack_8_wvalid & _writeStack_entryFifoid_T_51 & _canAW_T_50; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_53 = writeStack_8_wvalid & _writeStack_entryFifoid_T_51 & _canAW_T_50 & _canAW_T_52; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_57 = writeStack_9_wvalid & _writeStack_entryFifoid_T_57 & _canAW_T_56; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_59 = writeStack_9_wvalid & _writeStack_entryFifoid_T_57 & _canAW_T_56 & _canAW_T_58; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_63 = writeStack_10_wvalid & _writeStack_entryFifoid_T_63 & _canAW_T_62; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_65 = writeStack_10_wvalid & _writeStack_entryFifoid_T_63 & _canAW_T_62 & _canAW_T_64; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_69 = writeStack_11_wvalid & _writeStack_entryFifoid_T_69 & _canAW_T_68; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_71 = writeStack_11_wvalid & _writeStack_entryFifoid_T_69 & _canAW_T_68 & _canAW_T_70; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_75 = writeStack_12_wvalid & _writeStack_entryFifoid_T_75 & _canAW_T_74; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_77 = writeStack_12_wvalid & _writeStack_entryFifoid_T_75 & _canAW_T_74 & _canAW_T_76; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_81 = writeStack_13_wvalid & _writeStack_entryFifoid_T_81 & _canAW_T_80; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_83 = writeStack_13_wvalid & _writeStack_entryFifoid_T_81 & _canAW_T_80 & _canAW_T_82; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_87 = writeStack_14_wvalid & _writeStack_entryFifoid_T_87 & _canAW_T_86; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_89 = writeStack_14_wvalid & _writeStack_entryFifoid_T_87 & _canAW_T_86 & _canAW_T_88; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_93 = writeStack_15_wvalid & _writeStack_entryFifoid_T_93 & _canAW_T_92; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_95 = writeStack_15_wvalid & _writeStack_entryFifoid_T_93 & _canAW_T_92 & _canAW_T_94; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_99 = writeStack_16_wvalid & _writeStack_entryFifoid_T_99 & _canAW_T_98; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_101 = writeStack_16_wvalid & _writeStack_entryFifoid_T_99 & _canAW_T_98 & _canAW_T_100; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_105 = writeStack_17_wvalid & _writeStack_entryFifoid_T_105 & _canAW_T_104; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_107 = writeStack_17_wvalid & _writeStack_entryFifoid_T_105 & _canAW_T_104 & _canAW_T_106; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_111 = writeStack_18_wvalid & _writeStack_entryFifoid_T_111 & _canAW_T_110; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_113 = writeStack_18_wvalid & _writeStack_entryFifoid_T_111 & _canAW_T_110 & _canAW_T_112; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_117 = writeStack_19_wvalid & _writeStack_entryFifoid_T_117 & _canAW_T_116; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_119 = writeStack_19_wvalid & _writeStack_entryFifoid_T_117 & _canAW_T_116 & _canAW_T_118; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_123 = writeStack_20_wvalid & _writeStack_entryFifoid_T_123 & _canAW_T_122; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_125 = writeStack_20_wvalid & _writeStack_entryFifoid_T_123 & _canAW_T_122 & _canAW_T_124; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_129 = writeStack_21_wvalid & _writeStack_entryFifoid_T_129 & _canAW_T_128; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_131 = writeStack_21_wvalid & _writeStack_entryFifoid_T_129 & _canAW_T_128 & _canAW_T_130; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_135 = writeStack_22_wvalid & _writeStack_entryFifoid_T_135 & _canAW_T_134; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_137 = writeStack_22_wvalid & _writeStack_entryFifoid_T_135 & _canAW_T_134 & _canAW_T_136; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_141 = writeStack_23_wvalid & _writeStack_entryFifoid_T_141 & _canAW_T_140; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_143 = writeStack_23_wvalid & _writeStack_entryFifoid_T_141 & _canAW_T_140 & _canAW_T_142; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_147 = writeStack_24_wvalid & _writeStack_entryFifoid_T_147 & _canAW_T_146; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_149 = writeStack_24_wvalid & _writeStack_entryFifoid_T_147 & _canAW_T_146 & _canAW_T_148; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_153 = writeStack_25_wvalid & _writeStack_entryFifoid_T_153 & _canAW_T_152; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_155 = writeStack_25_wvalid & _writeStack_entryFifoid_T_153 & _canAW_T_152 & _canAW_T_154; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_159 = writeStack_26_wvalid & _writeStack_entryFifoid_T_159 & _canAW_T_158; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_161 = writeStack_26_wvalid & _writeStack_entryFifoid_T_159 & _canAW_T_158 & _canAW_T_160; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_165 = writeStack_27_wvalid & _writeStack_entryFifoid_T_165 & _canAW_T_164; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_167 = writeStack_27_wvalid & _writeStack_entryFifoid_T_165 & _canAW_T_164 & _canAW_T_166; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_171 = writeStack_28_wvalid & _writeStack_entryFifoid_T_171 & _canAW_T_170; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_173 = writeStack_28_wvalid & _writeStack_entryFifoid_T_171 & _canAW_T_170 & _canAW_T_172; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_177 = writeStack_29_wvalid & _writeStack_entryFifoid_T_177 & _canAW_T_176; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_179 = writeStack_29_wvalid & _writeStack_entryFifoid_T_177 & _canAW_T_176 & _canAW_T_178; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_183 = writeStack_30_wvalid & _writeStack_entryFifoid_T_183 & _canAW_T_182; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_185 = writeStack_30_wvalid & _writeStack_entryFifoid_T_183 & _canAW_T_182 & _canAW_T_184; // @[WriteStack.scala 213:104]
  wire  _canMenW_T_189 = writeStack_31_wvalid & _writeStack_entryFifoid_T_189 & _canAW_T_188; // @[WriteStack.scala 213:73]
  wire  _canMenW_T_191 = writeStack_31_wvalid & _writeStack_entryFifoid_T_189 & _canAW_T_188 & _canAW_T_190; // @[WriteStack.scala 213:104]
  wire [4:0] _writeStack_0_entryFifoid_T_1 = writeStack_0_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_609 = writeStack_0_wvalid & writeStack_0_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1537 = _canMenW_T_5 ? 3'h5 : _GEN_1504; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1539 = _canMenW_T_5 ? 3'h0 : {{1'd0}, _GEN_1312}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_1_entryFifoid_T_1 = writeStack_1_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_617 = writeStack_1_wvalid & writeStack_1_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1542 = _canMenW_T_11 ? 3'h5 : _GEN_1505; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1544 = _canMenW_T_11 ? 3'h0 : {{1'd0}, _GEN_1313}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_2_entryFifoid_T_1 = writeStack_2_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_625 = writeStack_2_wvalid & writeStack_2_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1547 = _canMenW_T_17 ? 3'h5 : _GEN_1506; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1549 = _canMenW_T_17 ? 3'h0 : {{1'd0}, _GEN_1314}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_3_entryFifoid_T_1 = writeStack_3_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_633 = writeStack_3_wvalid & writeStack_3_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1552 = _canMenW_T_23 ? 3'h5 : _GEN_1507; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1554 = _canMenW_T_23 ? 3'h0 : {{1'd0}, _GEN_1315}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_4_entryFifoid_T_1 = writeStack_4_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_641 = writeStack_4_wvalid & writeStack_4_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1557 = _canMenW_T_29 ? 3'h5 : _GEN_1508; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1559 = _canMenW_T_29 ? 3'h0 : {{1'd0}, _GEN_1316}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_5_entryFifoid_T_1 = writeStack_5_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_649 = writeStack_5_wvalid & writeStack_5_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1562 = _canMenW_T_35 ? 3'h5 : _GEN_1509; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1564 = _canMenW_T_35 ? 3'h0 : {{1'd0}, _GEN_1317}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_6_entryFifoid_T_1 = writeStack_6_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_657 = writeStack_6_wvalid & writeStack_6_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1567 = _canMenW_T_41 ? 3'h5 : _GEN_1510; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1569 = _canMenW_T_41 ? 3'h0 : {{1'd0}, _GEN_1318}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_7_entryFifoid_T_1 = writeStack_7_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_665 = writeStack_7_wvalid & writeStack_7_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1572 = _canMenW_T_47 ? 3'h5 : _GEN_1511; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1574 = _canMenW_T_47 ? 3'h0 : {{1'd0}, _GEN_1319}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_8_entryFifoid_T_1 = writeStack_8_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_673 = writeStack_8_wvalid & writeStack_8_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1577 = _canMenW_T_53 ? 3'h5 : _GEN_1512; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1579 = _canMenW_T_53 ? 3'h0 : {{1'd0}, _GEN_1320}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_9_entryFifoid_T_1 = writeStack_9_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_681 = writeStack_9_wvalid & writeStack_9_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1582 = _canMenW_T_59 ? 3'h5 : _GEN_1513; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1584 = _canMenW_T_59 ? 3'h0 : {{1'd0}, _GEN_1321}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_10_entryFifoid_T_1 = writeStack_10_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_689 = writeStack_10_wvalid & writeStack_10_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1587 = _canMenW_T_65 ? 3'h5 : _GEN_1514; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1589 = _canMenW_T_65 ? 3'h0 : {{1'd0}, _GEN_1322}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_11_entryFifoid_T_1 = writeStack_11_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_697 = writeStack_11_wvalid & writeStack_11_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1592 = _canMenW_T_71 ? 3'h5 : _GEN_1515; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1594 = _canMenW_T_71 ? 3'h0 : {{1'd0}, _GEN_1323}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_12_entryFifoid_T_1 = writeStack_12_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_705 = writeStack_12_wvalid & writeStack_12_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1597 = _canMenW_T_77 ? 3'h5 : _GEN_1516; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1599 = _canMenW_T_77 ? 3'h0 : {{1'd0}, _GEN_1324}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_13_entryFifoid_T_1 = writeStack_13_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_713 = writeStack_13_wvalid & writeStack_13_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1602 = _canMenW_T_83 ? 3'h5 : _GEN_1517; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1604 = _canMenW_T_83 ? 3'h0 : {{1'd0}, _GEN_1325}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_14_entryFifoid_T_1 = writeStack_14_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_721 = writeStack_14_wvalid & writeStack_14_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1607 = _canMenW_T_89 ? 3'h5 : _GEN_1518; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1609 = _canMenW_T_89 ? 3'h0 : {{1'd0}, _GEN_1326}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_15_entryFifoid_T_1 = writeStack_15_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_729 = writeStack_15_wvalid & writeStack_15_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1612 = _canMenW_T_95 ? 3'h5 : _GEN_1519; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1614 = _canMenW_T_95 ? 3'h0 : {{1'd0}, _GEN_1327}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_16_entryFifoid_T_1 = writeStack_16_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_737 = writeStack_16_wvalid & writeStack_16_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1617 = _canMenW_T_101 ? 3'h5 : _GEN_1520; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1619 = _canMenW_T_101 ? 3'h0 : {{1'd0}, _GEN_1328}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_17_entryFifoid_T_1 = writeStack_17_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_745 = writeStack_17_wvalid & writeStack_17_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1622 = _canMenW_T_107 ? 3'h5 : _GEN_1521; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1624 = _canMenW_T_107 ? 3'h0 : {{1'd0}, _GEN_1329}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_18_entryFifoid_T_1 = writeStack_18_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_753 = writeStack_18_wvalid & writeStack_18_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1627 = _canMenW_T_113 ? 3'h5 : _GEN_1522; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1629 = _canMenW_T_113 ? 3'h0 : {{1'd0}, _GEN_1330}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_19_entryFifoid_T_1 = writeStack_19_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_761 = writeStack_19_wvalid & writeStack_19_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1632 = _canMenW_T_119 ? 3'h5 : _GEN_1523; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1634 = _canMenW_T_119 ? 3'h0 : {{1'd0}, _GEN_1331}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_20_entryFifoid_T_1 = writeStack_20_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_769 = writeStack_20_wvalid & writeStack_20_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1637 = _canMenW_T_125 ? 3'h5 : _GEN_1524; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1639 = _canMenW_T_125 ? 3'h0 : {{1'd0}, _GEN_1332}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_21_entryFifoid_T_1 = writeStack_21_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_777 = writeStack_21_wvalid & writeStack_21_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1642 = _canMenW_T_131 ? 3'h5 : _GEN_1525; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1644 = _canMenW_T_131 ? 3'h0 : {{1'd0}, _GEN_1333}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_22_entryFifoid_T_1 = writeStack_22_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_785 = writeStack_22_wvalid & writeStack_22_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1647 = _canMenW_T_137 ? 3'h5 : _GEN_1526; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1649 = _canMenW_T_137 ? 3'h0 : {{1'd0}, _GEN_1334}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_23_entryFifoid_T_1 = writeStack_23_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_793 = writeStack_23_wvalid & writeStack_23_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1652 = _canMenW_T_143 ? 3'h5 : _GEN_1527; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1654 = _canMenW_T_143 ? 3'h0 : {{1'd0}, _GEN_1335}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_24_entryFifoid_T_1 = writeStack_24_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_801 = writeStack_24_wvalid & writeStack_24_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1657 = _canMenW_T_149 ? 3'h5 : _GEN_1528; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1659 = _canMenW_T_149 ? 3'h0 : {{1'd0}, _GEN_1336}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_25_entryFifoid_T_1 = writeStack_25_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_809 = writeStack_25_wvalid & writeStack_25_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1662 = _canMenW_T_155 ? 3'h5 : _GEN_1529; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1664 = _canMenW_T_155 ? 3'h0 : {{1'd0}, _GEN_1337}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_26_entryFifoid_T_1 = writeStack_26_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_817 = writeStack_26_wvalid & writeStack_26_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1667 = _canMenW_T_161 ? 3'h5 : _GEN_1530; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1669 = _canMenW_T_161 ? 3'h0 : {{1'd0}, _GEN_1338}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_27_entryFifoid_T_1 = writeStack_27_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_825 = writeStack_27_wvalid & writeStack_27_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1672 = _canMenW_T_167 ? 3'h5 : _GEN_1531; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1674 = _canMenW_T_167 ? 3'h0 : {{1'd0}, _GEN_1339}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_28_entryFifoid_T_1 = writeStack_28_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_833 = writeStack_28_wvalid & writeStack_28_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1677 = _canMenW_T_173 ? 3'h5 : _GEN_1532; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1679 = _canMenW_T_173 ? 3'h0 : {{1'd0}, _GEN_1340}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_29_entryFifoid_T_1 = writeStack_29_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_841 = writeStack_29_wvalid & writeStack_29_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1682 = _canMenW_T_179 ? 3'h5 : _GEN_1533; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1684 = _canMenW_T_179 ? 3'h0 : {{1'd0}, _GEN_1341}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_30_entryFifoid_T_1 = writeStack_30_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_849 = writeStack_30_wvalid & writeStack_30_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1687 = _canMenW_T_185 ? 3'h5 : _GEN_1534; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1689 = _canMenW_T_185 ? 3'h0 : {{1'd0}, _GEN_1342}; // @[WriteStack.scala 233:15 237:33]
  wire [4:0] _writeStack_31_entryFifoid_T_1 = writeStack_31_entryFifoid - 5'h1; // @[WriteStack.scala 238:50]
  wire  _T_857 = writeStack_31_wvalid & writeStack_31_entryFifoid != 5'h0; // @[WriteStack.scala 239:36]
  wire [2:0] _GEN_1692 = _canMenW_T_191 ? 3'h5 : _GEN_1535; // @[WriteStack.scala 233:15 235:29]
  wire [2:0] _GEN_1694 = _canMenW_T_191 ? 3'h0 : {{1'd0}, _GEN_1343}; // @[WriteStack.scala 233:15 237:33]
  wire [2:0] _GEN_1696 = _T_402 ? _GEN_1537 : _GEN_1504; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1698 = _T_402 ? _GEN_1539 : {{1'd0}, _GEN_1312}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1700 = _T_402 ? _GEN_1542 : _GEN_1505; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1702 = _T_402 ? _GEN_1544 : {{1'd0}, _GEN_1313}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1704 = _T_402 ? _GEN_1547 : _GEN_1506; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1706 = _T_402 ? _GEN_1549 : {{1'd0}, _GEN_1314}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1708 = _T_402 ? _GEN_1552 : _GEN_1507; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1710 = _T_402 ? _GEN_1554 : {{1'd0}, _GEN_1315}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1712 = _T_402 ? _GEN_1557 : _GEN_1508; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1714 = _T_402 ? _GEN_1559 : {{1'd0}, _GEN_1316}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1716 = _T_402 ? _GEN_1562 : _GEN_1509; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1718 = _T_402 ? _GEN_1564 : {{1'd0}, _GEN_1317}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1720 = _T_402 ? _GEN_1567 : _GEN_1510; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1722 = _T_402 ? _GEN_1569 : {{1'd0}, _GEN_1318}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1724 = _T_402 ? _GEN_1572 : _GEN_1511; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1726 = _T_402 ? _GEN_1574 : {{1'd0}, _GEN_1319}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1728 = _T_402 ? _GEN_1577 : _GEN_1512; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1730 = _T_402 ? _GEN_1579 : {{1'd0}, _GEN_1320}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1732 = _T_402 ? _GEN_1582 : _GEN_1513; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1734 = _T_402 ? _GEN_1584 : {{1'd0}, _GEN_1321}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1736 = _T_402 ? _GEN_1587 : _GEN_1514; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1738 = _T_402 ? _GEN_1589 : {{1'd0}, _GEN_1322}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1740 = _T_402 ? _GEN_1592 : _GEN_1515; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1742 = _T_402 ? _GEN_1594 : {{1'd0}, _GEN_1323}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1744 = _T_402 ? _GEN_1597 : _GEN_1516; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1746 = _T_402 ? _GEN_1599 : {{1'd0}, _GEN_1324}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1748 = _T_402 ? _GEN_1602 : _GEN_1517; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1750 = _T_402 ? _GEN_1604 : {{1'd0}, _GEN_1325}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1752 = _T_402 ? _GEN_1607 : _GEN_1518; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1754 = _T_402 ? _GEN_1609 : {{1'd0}, _GEN_1326}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1756 = _T_402 ? _GEN_1612 : _GEN_1519; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1758 = _T_402 ? _GEN_1614 : {{1'd0}, _GEN_1327}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1760 = _T_402 ? _GEN_1617 : _GEN_1520; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1762 = _T_402 ? _GEN_1619 : {{1'd0}, _GEN_1328}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1764 = _T_402 ? _GEN_1622 : _GEN_1521; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1766 = _T_402 ? _GEN_1624 : {{1'd0}, _GEN_1329}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1768 = _T_402 ? _GEN_1627 : _GEN_1522; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1770 = _T_402 ? _GEN_1629 : {{1'd0}, _GEN_1330}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1772 = _T_402 ? _GEN_1632 : _GEN_1523; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1774 = _T_402 ? _GEN_1634 : {{1'd0}, _GEN_1331}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1776 = _T_402 ? _GEN_1637 : _GEN_1524; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1778 = _T_402 ? _GEN_1639 : {{1'd0}, _GEN_1332}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1780 = _T_402 ? _GEN_1642 : _GEN_1525; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1782 = _T_402 ? _GEN_1644 : {{1'd0}, _GEN_1333}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1784 = _T_402 ? _GEN_1647 : _GEN_1526; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1786 = _T_402 ? _GEN_1649 : {{1'd0}, _GEN_1334}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1788 = _T_402 ? _GEN_1652 : _GEN_1527; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1790 = _T_402 ? _GEN_1654 : {{1'd0}, _GEN_1335}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1792 = _T_402 ? _GEN_1657 : _GEN_1528; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1794 = _T_402 ? _GEN_1659 : {{1'd0}, _GEN_1336}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1796 = _T_402 ? _GEN_1662 : _GEN_1529; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1798 = _T_402 ? _GEN_1664 : {{1'd0}, _GEN_1337}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1800 = _T_402 ? _GEN_1667 : _GEN_1530; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1802 = _T_402 ? _GEN_1669 : {{1'd0}, _GEN_1338}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1804 = _T_402 ? _GEN_1672 : _GEN_1531; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1806 = _T_402 ? _GEN_1674 : {{1'd0}, _GEN_1339}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1808 = _T_402 ? _GEN_1677 : _GEN_1532; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1810 = _T_402 ? _GEN_1679 : {{1'd0}, _GEN_1340}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1812 = _T_402 ? _GEN_1682 : _GEN_1533; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1814 = _T_402 ? _GEN_1684 : {{1'd0}, _GEN_1341}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1816 = _T_402 ? _GEN_1687 : _GEN_1534; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1818 = _T_402 ? _GEN_1689 : {{1'd0}, _GEN_1342}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1820 = _T_402 ? _GEN_1692 : _GEN_1535; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_1822 = _T_402 ? _GEN_1694 : {{1'd0}, _GEN_1343}; // @[WriteStack.scala 229:3]
  wire [2:0] _GEN_2432 = reset ? 3'h0 : _GEN_1696; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2433 = reset ? 3'h0 : _GEN_1698; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2434 = reset ? 3'h0 : _GEN_1700; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2435 = reset ? 3'h0 : _GEN_1702; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2436 = reset ? 3'h0 : _GEN_1704; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2437 = reset ? 3'h0 : _GEN_1706; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2438 = reset ? 3'h0 : _GEN_1708; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2439 = reset ? 3'h0 : _GEN_1710; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2440 = reset ? 3'h0 : _GEN_1712; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2441 = reset ? 3'h0 : _GEN_1714; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2442 = reset ? 3'h0 : _GEN_1716; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2443 = reset ? 3'h0 : _GEN_1718; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2444 = reset ? 3'h0 : _GEN_1720; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2445 = reset ? 3'h0 : _GEN_1722; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2446 = reset ? 3'h0 : _GEN_1724; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2447 = reset ? 3'h0 : _GEN_1726; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2448 = reset ? 3'h0 : _GEN_1728; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2449 = reset ? 3'h0 : _GEN_1730; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2450 = reset ? 3'h0 : _GEN_1732; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2451 = reset ? 3'h0 : _GEN_1734; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2452 = reset ? 3'h0 : _GEN_1736; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2453 = reset ? 3'h0 : _GEN_1738; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2454 = reset ? 3'h0 : _GEN_1740; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2455 = reset ? 3'h0 : _GEN_1742; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2456 = reset ? 3'h0 : _GEN_1744; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2457 = reset ? 3'h0 : _GEN_1746; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2458 = reset ? 3'h0 : _GEN_1748; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2459 = reset ? 3'h0 : _GEN_1750; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2460 = reset ? 3'h0 : _GEN_1752; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2461 = reset ? 3'h0 : _GEN_1754; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2462 = reset ? 3'h0 : _GEN_1756; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2463 = reset ? 3'h0 : _GEN_1758; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2464 = reset ? 3'h0 : _GEN_1760; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2465 = reset ? 3'h0 : _GEN_1762; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2466 = reset ? 3'h0 : _GEN_1764; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2467 = reset ? 3'h0 : _GEN_1766; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2468 = reset ? 3'h0 : _GEN_1768; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2469 = reset ? 3'h0 : _GEN_1770; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2470 = reset ? 3'h0 : _GEN_1772; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2471 = reset ? 3'h0 : _GEN_1774; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2472 = reset ? 3'h0 : _GEN_1776; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2473 = reset ? 3'h0 : _GEN_1778; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2474 = reset ? 3'h0 : _GEN_1780; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2475 = reset ? 3'h0 : _GEN_1782; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2476 = reset ? 3'h0 : _GEN_1784; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2477 = reset ? 3'h0 : _GEN_1786; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2478 = reset ? 3'h0 : _GEN_1788; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2479 = reset ? 3'h0 : _GEN_1790; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2480 = reset ? 3'h0 : _GEN_1792; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2481 = reset ? 3'h0 : _GEN_1794; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2482 = reset ? 3'h0 : _GEN_1796; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2483 = reset ? 3'h0 : _GEN_1798; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2484 = reset ? 3'h0 : _GEN_1800; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2485 = reset ? 3'h0 : _GEN_1802; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2486 = reset ? 3'h0 : _GEN_1804; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2487 = reset ? 3'h0 : _GEN_1806; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2488 = reset ? 3'h0 : _GEN_1808; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2489 = reset ? 3'h0 : _GEN_1810; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2490 = reset ? 3'h0 : _GEN_1812; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2491 = reset ? 3'h0 : _GEN_1814; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2492 = reset ? 3'h0 : _GEN_1816; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2493 = reset ? 3'h0 : _GEN_1818; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2494 = reset ? 3'h0 : _GEN_1820; // @[WriteStack.scala 56:{27,27}]
  wire [2:0] _GEN_2495 = reset ? 3'h0 : _GEN_1822; // @[WriteStack.scala 56:{27,27}]
  Arbiter wreqArb ( // @[WriteStack.scala 60:23]
    .io_in_0_valid(wreqArb_io_in_0_valid),
    .io_in_0_bits_waddr(wreqArb_io_in_0_bits_waddr),
    .io_in_0_bits_entryid(wreqArb_io_in_0_bits_entryid),
    .io_in_0_bits_awid(wreqArb_io_in_0_bits_awid),
    .io_in_0_bits_data(wreqArb_io_in_0_bits_data),
    .io_in_0_bits_mask(wreqArb_io_in_0_bits_mask),
    .io_in_0_bits_size(wreqArb_io_in_0_bits_size),
    .io_in_0_bits_len(wreqArb_io_in_0_bits_len),
    .io_in_1_valid(wreqArb_io_in_1_valid),
    .io_in_1_bits_waddr(wreqArb_io_in_1_bits_waddr),
    .io_in_1_bits_entryid(wreqArb_io_in_1_bits_entryid),
    .io_in_1_bits_awid(wreqArb_io_in_1_bits_awid),
    .io_in_1_bits_data(wreqArb_io_in_1_bits_data),
    .io_in_1_bits_mask(wreqArb_io_in_1_bits_mask),
    .io_in_1_bits_size(wreqArb_io_in_1_bits_size),
    .io_in_1_bits_len(wreqArb_io_in_1_bits_len),
    .io_in_2_valid(wreqArb_io_in_2_valid),
    .io_in_2_bits_waddr(wreqArb_io_in_2_bits_waddr),
    .io_in_2_bits_entryid(wreqArb_io_in_2_bits_entryid),
    .io_in_2_bits_awid(wreqArb_io_in_2_bits_awid),
    .io_in_2_bits_data(wreqArb_io_in_2_bits_data),
    .io_in_2_bits_mask(wreqArb_io_in_2_bits_mask),
    .io_in_2_bits_size(wreqArb_io_in_2_bits_size),
    .io_in_2_bits_len(wreqArb_io_in_2_bits_len),
    .io_in_3_valid(wreqArb_io_in_3_valid),
    .io_in_3_bits_waddr(wreqArb_io_in_3_bits_waddr),
    .io_in_3_bits_entryid(wreqArb_io_in_3_bits_entryid),
    .io_in_3_bits_awid(wreqArb_io_in_3_bits_awid),
    .io_in_3_bits_data(wreqArb_io_in_3_bits_data),
    .io_in_3_bits_mask(wreqArb_io_in_3_bits_mask),
    .io_in_3_bits_size(wreqArb_io_in_3_bits_size),
    .io_in_3_bits_len(wreqArb_io_in_3_bits_len),
    .io_in_4_valid(wreqArb_io_in_4_valid),
    .io_in_4_bits_waddr(wreqArb_io_in_4_bits_waddr),
    .io_in_4_bits_entryid(wreqArb_io_in_4_bits_entryid),
    .io_in_4_bits_awid(wreqArb_io_in_4_bits_awid),
    .io_in_4_bits_data(wreqArb_io_in_4_bits_data),
    .io_in_4_bits_mask(wreqArb_io_in_4_bits_mask),
    .io_in_4_bits_size(wreqArb_io_in_4_bits_size),
    .io_in_4_bits_len(wreqArb_io_in_4_bits_len),
    .io_in_5_valid(wreqArb_io_in_5_valid),
    .io_in_5_bits_waddr(wreqArb_io_in_5_bits_waddr),
    .io_in_5_bits_entryid(wreqArb_io_in_5_bits_entryid),
    .io_in_5_bits_awid(wreqArb_io_in_5_bits_awid),
    .io_in_5_bits_data(wreqArb_io_in_5_bits_data),
    .io_in_5_bits_mask(wreqArb_io_in_5_bits_mask),
    .io_in_5_bits_size(wreqArb_io_in_5_bits_size),
    .io_in_5_bits_len(wreqArb_io_in_5_bits_len),
    .io_in_6_valid(wreqArb_io_in_6_valid),
    .io_in_6_bits_waddr(wreqArb_io_in_6_bits_waddr),
    .io_in_6_bits_entryid(wreqArb_io_in_6_bits_entryid),
    .io_in_6_bits_awid(wreqArb_io_in_6_bits_awid),
    .io_in_6_bits_data(wreqArb_io_in_6_bits_data),
    .io_in_6_bits_mask(wreqArb_io_in_6_bits_mask),
    .io_in_6_bits_size(wreqArb_io_in_6_bits_size),
    .io_in_6_bits_len(wreqArb_io_in_6_bits_len),
    .io_in_7_valid(wreqArb_io_in_7_valid),
    .io_in_7_bits_waddr(wreqArb_io_in_7_bits_waddr),
    .io_in_7_bits_entryid(wreqArb_io_in_7_bits_entryid),
    .io_in_7_bits_awid(wreqArb_io_in_7_bits_awid),
    .io_in_7_bits_data(wreqArb_io_in_7_bits_data),
    .io_in_7_bits_mask(wreqArb_io_in_7_bits_mask),
    .io_in_7_bits_size(wreqArb_io_in_7_bits_size),
    .io_in_7_bits_len(wreqArb_io_in_7_bits_len),
    .io_in_8_valid(wreqArb_io_in_8_valid),
    .io_in_8_bits_waddr(wreqArb_io_in_8_bits_waddr),
    .io_in_8_bits_entryid(wreqArb_io_in_8_bits_entryid),
    .io_in_8_bits_awid(wreqArb_io_in_8_bits_awid),
    .io_in_8_bits_data(wreqArb_io_in_8_bits_data),
    .io_in_8_bits_mask(wreqArb_io_in_8_bits_mask),
    .io_in_8_bits_size(wreqArb_io_in_8_bits_size),
    .io_in_8_bits_len(wreqArb_io_in_8_bits_len),
    .io_in_9_valid(wreqArb_io_in_9_valid),
    .io_in_9_bits_waddr(wreqArb_io_in_9_bits_waddr),
    .io_in_9_bits_entryid(wreqArb_io_in_9_bits_entryid),
    .io_in_9_bits_awid(wreqArb_io_in_9_bits_awid),
    .io_in_9_bits_data(wreqArb_io_in_9_bits_data),
    .io_in_9_bits_mask(wreqArb_io_in_9_bits_mask),
    .io_in_9_bits_size(wreqArb_io_in_9_bits_size),
    .io_in_9_bits_len(wreqArb_io_in_9_bits_len),
    .io_in_10_valid(wreqArb_io_in_10_valid),
    .io_in_10_bits_waddr(wreqArb_io_in_10_bits_waddr),
    .io_in_10_bits_entryid(wreqArb_io_in_10_bits_entryid),
    .io_in_10_bits_awid(wreqArb_io_in_10_bits_awid),
    .io_in_10_bits_data(wreqArb_io_in_10_bits_data),
    .io_in_10_bits_mask(wreqArb_io_in_10_bits_mask),
    .io_in_10_bits_size(wreqArb_io_in_10_bits_size),
    .io_in_10_bits_len(wreqArb_io_in_10_bits_len),
    .io_in_11_valid(wreqArb_io_in_11_valid),
    .io_in_11_bits_waddr(wreqArb_io_in_11_bits_waddr),
    .io_in_11_bits_entryid(wreqArb_io_in_11_bits_entryid),
    .io_in_11_bits_awid(wreqArb_io_in_11_bits_awid),
    .io_in_11_bits_data(wreqArb_io_in_11_bits_data),
    .io_in_11_bits_mask(wreqArb_io_in_11_bits_mask),
    .io_in_11_bits_size(wreqArb_io_in_11_bits_size),
    .io_in_11_bits_len(wreqArb_io_in_11_bits_len),
    .io_in_12_valid(wreqArb_io_in_12_valid),
    .io_in_12_bits_waddr(wreqArb_io_in_12_bits_waddr),
    .io_in_12_bits_entryid(wreqArb_io_in_12_bits_entryid),
    .io_in_12_bits_awid(wreqArb_io_in_12_bits_awid),
    .io_in_12_bits_data(wreqArb_io_in_12_bits_data),
    .io_in_12_bits_mask(wreqArb_io_in_12_bits_mask),
    .io_in_12_bits_size(wreqArb_io_in_12_bits_size),
    .io_in_12_bits_len(wreqArb_io_in_12_bits_len),
    .io_in_13_valid(wreqArb_io_in_13_valid),
    .io_in_13_bits_waddr(wreqArb_io_in_13_bits_waddr),
    .io_in_13_bits_entryid(wreqArb_io_in_13_bits_entryid),
    .io_in_13_bits_awid(wreqArb_io_in_13_bits_awid),
    .io_in_13_bits_data(wreqArb_io_in_13_bits_data),
    .io_in_13_bits_mask(wreqArb_io_in_13_bits_mask),
    .io_in_13_bits_size(wreqArb_io_in_13_bits_size),
    .io_in_13_bits_len(wreqArb_io_in_13_bits_len),
    .io_in_14_valid(wreqArb_io_in_14_valid),
    .io_in_14_bits_waddr(wreqArb_io_in_14_bits_waddr),
    .io_in_14_bits_entryid(wreqArb_io_in_14_bits_entryid),
    .io_in_14_bits_awid(wreqArb_io_in_14_bits_awid),
    .io_in_14_bits_data(wreqArb_io_in_14_bits_data),
    .io_in_14_bits_mask(wreqArb_io_in_14_bits_mask),
    .io_in_14_bits_size(wreqArb_io_in_14_bits_size),
    .io_in_14_bits_len(wreqArb_io_in_14_bits_len),
    .io_in_15_valid(wreqArb_io_in_15_valid),
    .io_in_15_bits_waddr(wreqArb_io_in_15_bits_waddr),
    .io_in_15_bits_entryid(wreqArb_io_in_15_bits_entryid),
    .io_in_15_bits_awid(wreqArb_io_in_15_bits_awid),
    .io_in_15_bits_data(wreqArb_io_in_15_bits_data),
    .io_in_15_bits_mask(wreqArb_io_in_15_bits_mask),
    .io_in_15_bits_size(wreqArb_io_in_15_bits_size),
    .io_in_15_bits_len(wreqArb_io_in_15_bits_len),
    .io_in_16_valid(wreqArb_io_in_16_valid),
    .io_in_16_bits_waddr(wreqArb_io_in_16_bits_waddr),
    .io_in_16_bits_entryid(wreqArb_io_in_16_bits_entryid),
    .io_in_16_bits_awid(wreqArb_io_in_16_bits_awid),
    .io_in_16_bits_data(wreqArb_io_in_16_bits_data),
    .io_in_16_bits_mask(wreqArb_io_in_16_bits_mask),
    .io_in_16_bits_size(wreqArb_io_in_16_bits_size),
    .io_in_16_bits_len(wreqArb_io_in_16_bits_len),
    .io_in_17_valid(wreqArb_io_in_17_valid),
    .io_in_17_bits_waddr(wreqArb_io_in_17_bits_waddr),
    .io_in_17_bits_entryid(wreqArb_io_in_17_bits_entryid),
    .io_in_17_bits_awid(wreqArb_io_in_17_bits_awid),
    .io_in_17_bits_data(wreqArb_io_in_17_bits_data),
    .io_in_17_bits_mask(wreqArb_io_in_17_bits_mask),
    .io_in_17_bits_size(wreqArb_io_in_17_bits_size),
    .io_in_17_bits_len(wreqArb_io_in_17_bits_len),
    .io_in_18_valid(wreqArb_io_in_18_valid),
    .io_in_18_bits_waddr(wreqArb_io_in_18_bits_waddr),
    .io_in_18_bits_entryid(wreqArb_io_in_18_bits_entryid),
    .io_in_18_bits_awid(wreqArb_io_in_18_bits_awid),
    .io_in_18_bits_data(wreqArb_io_in_18_bits_data),
    .io_in_18_bits_mask(wreqArb_io_in_18_bits_mask),
    .io_in_18_bits_size(wreqArb_io_in_18_bits_size),
    .io_in_18_bits_len(wreqArb_io_in_18_bits_len),
    .io_in_19_valid(wreqArb_io_in_19_valid),
    .io_in_19_bits_waddr(wreqArb_io_in_19_bits_waddr),
    .io_in_19_bits_entryid(wreqArb_io_in_19_bits_entryid),
    .io_in_19_bits_awid(wreqArb_io_in_19_bits_awid),
    .io_in_19_bits_data(wreqArb_io_in_19_bits_data),
    .io_in_19_bits_mask(wreqArb_io_in_19_bits_mask),
    .io_in_19_bits_size(wreqArb_io_in_19_bits_size),
    .io_in_19_bits_len(wreqArb_io_in_19_bits_len),
    .io_in_20_valid(wreqArb_io_in_20_valid),
    .io_in_20_bits_waddr(wreqArb_io_in_20_bits_waddr),
    .io_in_20_bits_entryid(wreqArb_io_in_20_bits_entryid),
    .io_in_20_bits_awid(wreqArb_io_in_20_bits_awid),
    .io_in_20_bits_data(wreqArb_io_in_20_bits_data),
    .io_in_20_bits_mask(wreqArb_io_in_20_bits_mask),
    .io_in_20_bits_size(wreqArb_io_in_20_bits_size),
    .io_in_20_bits_len(wreqArb_io_in_20_bits_len),
    .io_in_21_valid(wreqArb_io_in_21_valid),
    .io_in_21_bits_waddr(wreqArb_io_in_21_bits_waddr),
    .io_in_21_bits_entryid(wreqArb_io_in_21_bits_entryid),
    .io_in_21_bits_awid(wreqArb_io_in_21_bits_awid),
    .io_in_21_bits_data(wreqArb_io_in_21_bits_data),
    .io_in_21_bits_mask(wreqArb_io_in_21_bits_mask),
    .io_in_21_bits_size(wreqArb_io_in_21_bits_size),
    .io_in_21_bits_len(wreqArb_io_in_21_bits_len),
    .io_in_22_valid(wreqArb_io_in_22_valid),
    .io_in_22_bits_waddr(wreqArb_io_in_22_bits_waddr),
    .io_in_22_bits_entryid(wreqArb_io_in_22_bits_entryid),
    .io_in_22_bits_awid(wreqArb_io_in_22_bits_awid),
    .io_in_22_bits_data(wreqArb_io_in_22_bits_data),
    .io_in_22_bits_mask(wreqArb_io_in_22_bits_mask),
    .io_in_22_bits_size(wreqArb_io_in_22_bits_size),
    .io_in_22_bits_len(wreqArb_io_in_22_bits_len),
    .io_in_23_valid(wreqArb_io_in_23_valid),
    .io_in_23_bits_waddr(wreqArb_io_in_23_bits_waddr),
    .io_in_23_bits_entryid(wreqArb_io_in_23_bits_entryid),
    .io_in_23_bits_awid(wreqArb_io_in_23_bits_awid),
    .io_in_23_bits_data(wreqArb_io_in_23_bits_data),
    .io_in_23_bits_mask(wreqArb_io_in_23_bits_mask),
    .io_in_23_bits_size(wreqArb_io_in_23_bits_size),
    .io_in_23_bits_len(wreqArb_io_in_23_bits_len),
    .io_in_24_valid(wreqArb_io_in_24_valid),
    .io_in_24_bits_waddr(wreqArb_io_in_24_bits_waddr),
    .io_in_24_bits_entryid(wreqArb_io_in_24_bits_entryid),
    .io_in_24_bits_awid(wreqArb_io_in_24_bits_awid),
    .io_in_24_bits_data(wreqArb_io_in_24_bits_data),
    .io_in_24_bits_mask(wreqArb_io_in_24_bits_mask),
    .io_in_24_bits_size(wreqArb_io_in_24_bits_size),
    .io_in_24_bits_len(wreqArb_io_in_24_bits_len),
    .io_in_25_valid(wreqArb_io_in_25_valid),
    .io_in_25_bits_waddr(wreqArb_io_in_25_bits_waddr),
    .io_in_25_bits_entryid(wreqArb_io_in_25_bits_entryid),
    .io_in_25_bits_awid(wreqArb_io_in_25_bits_awid),
    .io_in_25_bits_data(wreqArb_io_in_25_bits_data),
    .io_in_25_bits_mask(wreqArb_io_in_25_bits_mask),
    .io_in_25_bits_size(wreqArb_io_in_25_bits_size),
    .io_in_25_bits_len(wreqArb_io_in_25_bits_len),
    .io_in_26_valid(wreqArb_io_in_26_valid),
    .io_in_26_bits_waddr(wreqArb_io_in_26_bits_waddr),
    .io_in_26_bits_entryid(wreqArb_io_in_26_bits_entryid),
    .io_in_26_bits_awid(wreqArb_io_in_26_bits_awid),
    .io_in_26_bits_data(wreqArb_io_in_26_bits_data),
    .io_in_26_bits_mask(wreqArb_io_in_26_bits_mask),
    .io_in_26_bits_size(wreqArb_io_in_26_bits_size),
    .io_in_26_bits_len(wreqArb_io_in_26_bits_len),
    .io_in_27_valid(wreqArb_io_in_27_valid),
    .io_in_27_bits_waddr(wreqArb_io_in_27_bits_waddr),
    .io_in_27_bits_entryid(wreqArb_io_in_27_bits_entryid),
    .io_in_27_bits_awid(wreqArb_io_in_27_bits_awid),
    .io_in_27_bits_data(wreqArb_io_in_27_bits_data),
    .io_in_27_bits_mask(wreqArb_io_in_27_bits_mask),
    .io_in_27_bits_size(wreqArb_io_in_27_bits_size),
    .io_in_27_bits_len(wreqArb_io_in_27_bits_len),
    .io_in_28_valid(wreqArb_io_in_28_valid),
    .io_in_28_bits_waddr(wreqArb_io_in_28_bits_waddr),
    .io_in_28_bits_entryid(wreqArb_io_in_28_bits_entryid),
    .io_in_28_bits_awid(wreqArb_io_in_28_bits_awid),
    .io_in_28_bits_data(wreqArb_io_in_28_bits_data),
    .io_in_28_bits_mask(wreqArb_io_in_28_bits_mask),
    .io_in_28_bits_size(wreqArb_io_in_28_bits_size),
    .io_in_28_bits_len(wreqArb_io_in_28_bits_len),
    .io_in_29_valid(wreqArb_io_in_29_valid),
    .io_in_29_bits_waddr(wreqArb_io_in_29_bits_waddr),
    .io_in_29_bits_entryid(wreqArb_io_in_29_bits_entryid),
    .io_in_29_bits_awid(wreqArb_io_in_29_bits_awid),
    .io_in_29_bits_data(wreqArb_io_in_29_bits_data),
    .io_in_29_bits_mask(wreqArb_io_in_29_bits_mask),
    .io_in_29_bits_size(wreqArb_io_in_29_bits_size),
    .io_in_29_bits_len(wreqArb_io_in_29_bits_len),
    .io_in_30_valid(wreqArb_io_in_30_valid),
    .io_in_30_bits_waddr(wreqArb_io_in_30_bits_waddr),
    .io_in_30_bits_entryid(wreqArb_io_in_30_bits_entryid),
    .io_in_30_bits_awid(wreqArb_io_in_30_bits_awid),
    .io_in_30_bits_data(wreqArb_io_in_30_bits_data),
    .io_in_30_bits_mask(wreqArb_io_in_30_bits_mask),
    .io_in_30_bits_size(wreqArb_io_in_30_bits_size),
    .io_in_30_bits_len(wreqArb_io_in_30_bits_len),
    .io_in_31_valid(wreqArb_io_in_31_valid),
    .io_in_31_bits_waddr(wreqArb_io_in_31_bits_waddr),
    .io_in_31_bits_entryid(wreqArb_io_in_31_bits_entryid),
    .io_in_31_bits_awid(wreqArb_io_in_31_bits_awid),
    .io_in_31_bits_data(wreqArb_io_in_31_bits_data),
    .io_in_31_bits_mask(wreqArb_io_in_31_bits_mask),
    .io_in_31_bits_size(wreqArb_io_in_31_bits_size),
    .io_in_31_bits_len(wreqArb_io_in_31_bits_len),
    .io_out_valid(wreqArb_io_out_valid),
    .io_out_bits_waddr(wreqArb_io_out_bits_waddr),
    .io_out_bits_entryid(wreqArb_io_out_bits_entryid),
    .io_out_bits_awid(wreqArb_io_out_bits_awid),
    .io_out_bits_data(wreqArb_io_out_bits_data),
    .io_out_bits_mask(wreqArb_io_out_bits_mask),
    .io_out_bits_size(wreqArb_io_out_bits_size),
    .io_out_bits_len(wreqArb_io_out_bits_len)
  );
  Arbiter awreqArb ( // @[WriteStack.scala 61:24]
    .io_in_0_valid(awreqArb_io_in_0_valid),
    .io_in_0_bits_waddr(awreqArb_io_in_0_bits_waddr),
    .io_in_0_bits_entryid(awreqArb_io_in_0_bits_entryid),
    .io_in_0_bits_awid(awreqArb_io_in_0_bits_awid),
    .io_in_0_bits_data(awreqArb_io_in_0_bits_data),
    .io_in_0_bits_mask(awreqArb_io_in_0_bits_mask),
    .io_in_0_bits_size(awreqArb_io_in_0_bits_size),
    .io_in_0_bits_len(awreqArb_io_in_0_bits_len),
    .io_in_1_valid(awreqArb_io_in_1_valid),
    .io_in_1_bits_waddr(awreqArb_io_in_1_bits_waddr),
    .io_in_1_bits_entryid(awreqArb_io_in_1_bits_entryid),
    .io_in_1_bits_awid(awreqArb_io_in_1_bits_awid),
    .io_in_1_bits_data(awreqArb_io_in_1_bits_data),
    .io_in_1_bits_mask(awreqArb_io_in_1_bits_mask),
    .io_in_1_bits_size(awreqArb_io_in_1_bits_size),
    .io_in_1_bits_len(awreqArb_io_in_1_bits_len),
    .io_in_2_valid(awreqArb_io_in_2_valid),
    .io_in_2_bits_waddr(awreqArb_io_in_2_bits_waddr),
    .io_in_2_bits_entryid(awreqArb_io_in_2_bits_entryid),
    .io_in_2_bits_awid(awreqArb_io_in_2_bits_awid),
    .io_in_2_bits_data(awreqArb_io_in_2_bits_data),
    .io_in_2_bits_mask(awreqArb_io_in_2_bits_mask),
    .io_in_2_bits_size(awreqArb_io_in_2_bits_size),
    .io_in_2_bits_len(awreqArb_io_in_2_bits_len),
    .io_in_3_valid(awreqArb_io_in_3_valid),
    .io_in_3_bits_waddr(awreqArb_io_in_3_bits_waddr),
    .io_in_3_bits_entryid(awreqArb_io_in_3_bits_entryid),
    .io_in_3_bits_awid(awreqArb_io_in_3_bits_awid),
    .io_in_3_bits_data(awreqArb_io_in_3_bits_data),
    .io_in_3_bits_mask(awreqArb_io_in_3_bits_mask),
    .io_in_3_bits_size(awreqArb_io_in_3_bits_size),
    .io_in_3_bits_len(awreqArb_io_in_3_bits_len),
    .io_in_4_valid(awreqArb_io_in_4_valid),
    .io_in_4_bits_waddr(awreqArb_io_in_4_bits_waddr),
    .io_in_4_bits_entryid(awreqArb_io_in_4_bits_entryid),
    .io_in_4_bits_awid(awreqArb_io_in_4_bits_awid),
    .io_in_4_bits_data(awreqArb_io_in_4_bits_data),
    .io_in_4_bits_mask(awreqArb_io_in_4_bits_mask),
    .io_in_4_bits_size(awreqArb_io_in_4_bits_size),
    .io_in_4_bits_len(awreqArb_io_in_4_bits_len),
    .io_in_5_valid(awreqArb_io_in_5_valid),
    .io_in_5_bits_waddr(awreqArb_io_in_5_bits_waddr),
    .io_in_5_bits_entryid(awreqArb_io_in_5_bits_entryid),
    .io_in_5_bits_awid(awreqArb_io_in_5_bits_awid),
    .io_in_5_bits_data(awreqArb_io_in_5_bits_data),
    .io_in_5_bits_mask(awreqArb_io_in_5_bits_mask),
    .io_in_5_bits_size(awreqArb_io_in_5_bits_size),
    .io_in_5_bits_len(awreqArb_io_in_5_bits_len),
    .io_in_6_valid(awreqArb_io_in_6_valid),
    .io_in_6_bits_waddr(awreqArb_io_in_6_bits_waddr),
    .io_in_6_bits_entryid(awreqArb_io_in_6_bits_entryid),
    .io_in_6_bits_awid(awreqArb_io_in_6_bits_awid),
    .io_in_6_bits_data(awreqArb_io_in_6_bits_data),
    .io_in_6_bits_mask(awreqArb_io_in_6_bits_mask),
    .io_in_6_bits_size(awreqArb_io_in_6_bits_size),
    .io_in_6_bits_len(awreqArb_io_in_6_bits_len),
    .io_in_7_valid(awreqArb_io_in_7_valid),
    .io_in_7_bits_waddr(awreqArb_io_in_7_bits_waddr),
    .io_in_7_bits_entryid(awreqArb_io_in_7_bits_entryid),
    .io_in_7_bits_awid(awreqArb_io_in_7_bits_awid),
    .io_in_7_bits_data(awreqArb_io_in_7_bits_data),
    .io_in_7_bits_mask(awreqArb_io_in_7_bits_mask),
    .io_in_7_bits_size(awreqArb_io_in_7_bits_size),
    .io_in_7_bits_len(awreqArb_io_in_7_bits_len),
    .io_in_8_valid(awreqArb_io_in_8_valid),
    .io_in_8_bits_waddr(awreqArb_io_in_8_bits_waddr),
    .io_in_8_bits_entryid(awreqArb_io_in_8_bits_entryid),
    .io_in_8_bits_awid(awreqArb_io_in_8_bits_awid),
    .io_in_8_bits_data(awreqArb_io_in_8_bits_data),
    .io_in_8_bits_mask(awreqArb_io_in_8_bits_mask),
    .io_in_8_bits_size(awreqArb_io_in_8_bits_size),
    .io_in_8_bits_len(awreqArb_io_in_8_bits_len),
    .io_in_9_valid(awreqArb_io_in_9_valid),
    .io_in_9_bits_waddr(awreqArb_io_in_9_bits_waddr),
    .io_in_9_bits_entryid(awreqArb_io_in_9_bits_entryid),
    .io_in_9_bits_awid(awreqArb_io_in_9_bits_awid),
    .io_in_9_bits_data(awreqArb_io_in_9_bits_data),
    .io_in_9_bits_mask(awreqArb_io_in_9_bits_mask),
    .io_in_9_bits_size(awreqArb_io_in_9_bits_size),
    .io_in_9_bits_len(awreqArb_io_in_9_bits_len),
    .io_in_10_valid(awreqArb_io_in_10_valid),
    .io_in_10_bits_waddr(awreqArb_io_in_10_bits_waddr),
    .io_in_10_bits_entryid(awreqArb_io_in_10_bits_entryid),
    .io_in_10_bits_awid(awreqArb_io_in_10_bits_awid),
    .io_in_10_bits_data(awreqArb_io_in_10_bits_data),
    .io_in_10_bits_mask(awreqArb_io_in_10_bits_mask),
    .io_in_10_bits_size(awreqArb_io_in_10_bits_size),
    .io_in_10_bits_len(awreqArb_io_in_10_bits_len),
    .io_in_11_valid(awreqArb_io_in_11_valid),
    .io_in_11_bits_waddr(awreqArb_io_in_11_bits_waddr),
    .io_in_11_bits_entryid(awreqArb_io_in_11_bits_entryid),
    .io_in_11_bits_awid(awreqArb_io_in_11_bits_awid),
    .io_in_11_bits_data(awreqArb_io_in_11_bits_data),
    .io_in_11_bits_mask(awreqArb_io_in_11_bits_mask),
    .io_in_11_bits_size(awreqArb_io_in_11_bits_size),
    .io_in_11_bits_len(awreqArb_io_in_11_bits_len),
    .io_in_12_valid(awreqArb_io_in_12_valid),
    .io_in_12_bits_waddr(awreqArb_io_in_12_bits_waddr),
    .io_in_12_bits_entryid(awreqArb_io_in_12_bits_entryid),
    .io_in_12_bits_awid(awreqArb_io_in_12_bits_awid),
    .io_in_12_bits_data(awreqArb_io_in_12_bits_data),
    .io_in_12_bits_mask(awreqArb_io_in_12_bits_mask),
    .io_in_12_bits_size(awreqArb_io_in_12_bits_size),
    .io_in_12_bits_len(awreqArb_io_in_12_bits_len),
    .io_in_13_valid(awreqArb_io_in_13_valid),
    .io_in_13_bits_waddr(awreqArb_io_in_13_bits_waddr),
    .io_in_13_bits_entryid(awreqArb_io_in_13_bits_entryid),
    .io_in_13_bits_awid(awreqArb_io_in_13_bits_awid),
    .io_in_13_bits_data(awreqArb_io_in_13_bits_data),
    .io_in_13_bits_mask(awreqArb_io_in_13_bits_mask),
    .io_in_13_bits_size(awreqArb_io_in_13_bits_size),
    .io_in_13_bits_len(awreqArb_io_in_13_bits_len),
    .io_in_14_valid(awreqArb_io_in_14_valid),
    .io_in_14_bits_waddr(awreqArb_io_in_14_bits_waddr),
    .io_in_14_bits_entryid(awreqArb_io_in_14_bits_entryid),
    .io_in_14_bits_awid(awreqArb_io_in_14_bits_awid),
    .io_in_14_bits_data(awreqArb_io_in_14_bits_data),
    .io_in_14_bits_mask(awreqArb_io_in_14_bits_mask),
    .io_in_14_bits_size(awreqArb_io_in_14_bits_size),
    .io_in_14_bits_len(awreqArb_io_in_14_bits_len),
    .io_in_15_valid(awreqArb_io_in_15_valid),
    .io_in_15_bits_waddr(awreqArb_io_in_15_bits_waddr),
    .io_in_15_bits_entryid(awreqArb_io_in_15_bits_entryid),
    .io_in_15_bits_awid(awreqArb_io_in_15_bits_awid),
    .io_in_15_bits_data(awreqArb_io_in_15_bits_data),
    .io_in_15_bits_mask(awreqArb_io_in_15_bits_mask),
    .io_in_15_bits_size(awreqArb_io_in_15_bits_size),
    .io_in_15_bits_len(awreqArb_io_in_15_bits_len),
    .io_in_16_valid(awreqArb_io_in_16_valid),
    .io_in_16_bits_waddr(awreqArb_io_in_16_bits_waddr),
    .io_in_16_bits_entryid(awreqArb_io_in_16_bits_entryid),
    .io_in_16_bits_awid(awreqArb_io_in_16_bits_awid),
    .io_in_16_bits_data(awreqArb_io_in_16_bits_data),
    .io_in_16_bits_mask(awreqArb_io_in_16_bits_mask),
    .io_in_16_bits_size(awreqArb_io_in_16_bits_size),
    .io_in_16_bits_len(awreqArb_io_in_16_bits_len),
    .io_in_17_valid(awreqArb_io_in_17_valid),
    .io_in_17_bits_waddr(awreqArb_io_in_17_bits_waddr),
    .io_in_17_bits_entryid(awreqArb_io_in_17_bits_entryid),
    .io_in_17_bits_awid(awreqArb_io_in_17_bits_awid),
    .io_in_17_bits_data(awreqArb_io_in_17_bits_data),
    .io_in_17_bits_mask(awreqArb_io_in_17_bits_mask),
    .io_in_17_bits_size(awreqArb_io_in_17_bits_size),
    .io_in_17_bits_len(awreqArb_io_in_17_bits_len),
    .io_in_18_valid(awreqArb_io_in_18_valid),
    .io_in_18_bits_waddr(awreqArb_io_in_18_bits_waddr),
    .io_in_18_bits_entryid(awreqArb_io_in_18_bits_entryid),
    .io_in_18_bits_awid(awreqArb_io_in_18_bits_awid),
    .io_in_18_bits_data(awreqArb_io_in_18_bits_data),
    .io_in_18_bits_mask(awreqArb_io_in_18_bits_mask),
    .io_in_18_bits_size(awreqArb_io_in_18_bits_size),
    .io_in_18_bits_len(awreqArb_io_in_18_bits_len),
    .io_in_19_valid(awreqArb_io_in_19_valid),
    .io_in_19_bits_waddr(awreqArb_io_in_19_bits_waddr),
    .io_in_19_bits_entryid(awreqArb_io_in_19_bits_entryid),
    .io_in_19_bits_awid(awreqArb_io_in_19_bits_awid),
    .io_in_19_bits_data(awreqArb_io_in_19_bits_data),
    .io_in_19_bits_mask(awreqArb_io_in_19_bits_mask),
    .io_in_19_bits_size(awreqArb_io_in_19_bits_size),
    .io_in_19_bits_len(awreqArb_io_in_19_bits_len),
    .io_in_20_valid(awreqArb_io_in_20_valid),
    .io_in_20_bits_waddr(awreqArb_io_in_20_bits_waddr),
    .io_in_20_bits_entryid(awreqArb_io_in_20_bits_entryid),
    .io_in_20_bits_awid(awreqArb_io_in_20_bits_awid),
    .io_in_20_bits_data(awreqArb_io_in_20_bits_data),
    .io_in_20_bits_mask(awreqArb_io_in_20_bits_mask),
    .io_in_20_bits_size(awreqArb_io_in_20_bits_size),
    .io_in_20_bits_len(awreqArb_io_in_20_bits_len),
    .io_in_21_valid(awreqArb_io_in_21_valid),
    .io_in_21_bits_waddr(awreqArb_io_in_21_bits_waddr),
    .io_in_21_bits_entryid(awreqArb_io_in_21_bits_entryid),
    .io_in_21_bits_awid(awreqArb_io_in_21_bits_awid),
    .io_in_21_bits_data(awreqArb_io_in_21_bits_data),
    .io_in_21_bits_mask(awreqArb_io_in_21_bits_mask),
    .io_in_21_bits_size(awreqArb_io_in_21_bits_size),
    .io_in_21_bits_len(awreqArb_io_in_21_bits_len),
    .io_in_22_valid(awreqArb_io_in_22_valid),
    .io_in_22_bits_waddr(awreqArb_io_in_22_bits_waddr),
    .io_in_22_bits_entryid(awreqArb_io_in_22_bits_entryid),
    .io_in_22_bits_awid(awreqArb_io_in_22_bits_awid),
    .io_in_22_bits_data(awreqArb_io_in_22_bits_data),
    .io_in_22_bits_mask(awreqArb_io_in_22_bits_mask),
    .io_in_22_bits_size(awreqArb_io_in_22_bits_size),
    .io_in_22_bits_len(awreqArb_io_in_22_bits_len),
    .io_in_23_valid(awreqArb_io_in_23_valid),
    .io_in_23_bits_waddr(awreqArb_io_in_23_bits_waddr),
    .io_in_23_bits_entryid(awreqArb_io_in_23_bits_entryid),
    .io_in_23_bits_awid(awreqArb_io_in_23_bits_awid),
    .io_in_23_bits_data(awreqArb_io_in_23_bits_data),
    .io_in_23_bits_mask(awreqArb_io_in_23_bits_mask),
    .io_in_23_bits_size(awreqArb_io_in_23_bits_size),
    .io_in_23_bits_len(awreqArb_io_in_23_bits_len),
    .io_in_24_valid(awreqArb_io_in_24_valid),
    .io_in_24_bits_waddr(awreqArb_io_in_24_bits_waddr),
    .io_in_24_bits_entryid(awreqArb_io_in_24_bits_entryid),
    .io_in_24_bits_awid(awreqArb_io_in_24_bits_awid),
    .io_in_24_bits_data(awreqArb_io_in_24_bits_data),
    .io_in_24_bits_mask(awreqArb_io_in_24_bits_mask),
    .io_in_24_bits_size(awreqArb_io_in_24_bits_size),
    .io_in_24_bits_len(awreqArb_io_in_24_bits_len),
    .io_in_25_valid(awreqArb_io_in_25_valid),
    .io_in_25_bits_waddr(awreqArb_io_in_25_bits_waddr),
    .io_in_25_bits_entryid(awreqArb_io_in_25_bits_entryid),
    .io_in_25_bits_awid(awreqArb_io_in_25_bits_awid),
    .io_in_25_bits_data(awreqArb_io_in_25_bits_data),
    .io_in_25_bits_mask(awreqArb_io_in_25_bits_mask),
    .io_in_25_bits_size(awreqArb_io_in_25_bits_size),
    .io_in_25_bits_len(awreqArb_io_in_25_bits_len),
    .io_in_26_valid(awreqArb_io_in_26_valid),
    .io_in_26_bits_waddr(awreqArb_io_in_26_bits_waddr),
    .io_in_26_bits_entryid(awreqArb_io_in_26_bits_entryid),
    .io_in_26_bits_awid(awreqArb_io_in_26_bits_awid),
    .io_in_26_bits_data(awreqArb_io_in_26_bits_data),
    .io_in_26_bits_mask(awreqArb_io_in_26_bits_mask),
    .io_in_26_bits_size(awreqArb_io_in_26_bits_size),
    .io_in_26_bits_len(awreqArb_io_in_26_bits_len),
    .io_in_27_valid(awreqArb_io_in_27_valid),
    .io_in_27_bits_waddr(awreqArb_io_in_27_bits_waddr),
    .io_in_27_bits_entryid(awreqArb_io_in_27_bits_entryid),
    .io_in_27_bits_awid(awreqArb_io_in_27_bits_awid),
    .io_in_27_bits_data(awreqArb_io_in_27_bits_data),
    .io_in_27_bits_mask(awreqArb_io_in_27_bits_mask),
    .io_in_27_bits_size(awreqArb_io_in_27_bits_size),
    .io_in_27_bits_len(awreqArb_io_in_27_bits_len),
    .io_in_28_valid(awreqArb_io_in_28_valid),
    .io_in_28_bits_waddr(awreqArb_io_in_28_bits_waddr),
    .io_in_28_bits_entryid(awreqArb_io_in_28_bits_entryid),
    .io_in_28_bits_awid(awreqArb_io_in_28_bits_awid),
    .io_in_28_bits_data(awreqArb_io_in_28_bits_data),
    .io_in_28_bits_mask(awreqArb_io_in_28_bits_mask),
    .io_in_28_bits_size(awreqArb_io_in_28_bits_size),
    .io_in_28_bits_len(awreqArb_io_in_28_bits_len),
    .io_in_29_valid(awreqArb_io_in_29_valid),
    .io_in_29_bits_waddr(awreqArb_io_in_29_bits_waddr),
    .io_in_29_bits_entryid(awreqArb_io_in_29_bits_entryid),
    .io_in_29_bits_awid(awreqArb_io_in_29_bits_awid),
    .io_in_29_bits_data(awreqArb_io_in_29_bits_data),
    .io_in_29_bits_mask(awreqArb_io_in_29_bits_mask),
    .io_in_29_bits_size(awreqArb_io_in_29_bits_size),
    .io_in_29_bits_len(awreqArb_io_in_29_bits_len),
    .io_in_30_valid(awreqArb_io_in_30_valid),
    .io_in_30_bits_waddr(awreqArb_io_in_30_bits_waddr),
    .io_in_30_bits_entryid(awreqArb_io_in_30_bits_entryid),
    .io_in_30_bits_awid(awreqArb_io_in_30_bits_awid),
    .io_in_30_bits_data(awreqArb_io_in_30_bits_data),
    .io_in_30_bits_mask(awreqArb_io_in_30_bits_mask),
    .io_in_30_bits_size(awreqArb_io_in_30_bits_size),
    .io_in_30_bits_len(awreqArb_io_in_30_bits_len),
    .io_in_31_valid(awreqArb_io_in_31_valid),
    .io_in_31_bits_waddr(awreqArb_io_in_31_bits_waddr),
    .io_in_31_bits_entryid(awreqArb_io_in_31_bits_entryid),
    .io_in_31_bits_awid(awreqArb_io_in_31_bits_awid),
    .io_in_31_bits_data(awreqArb_io_in_31_bits_data),
    .io_in_31_bits_mask(awreqArb_io_in_31_bits_mask),
    .io_in_31_bits_size(awreqArb_io_in_31_bits_size),
    .io_in_31_bits_len(awreqArb_io_in_31_bits_len),
    .io_out_valid(awreqArb_io_out_valid),
    .io_out_bits_waddr(awreqArb_io_out_bits_waddr),
    .io_out_bits_entryid(awreqArb_io_out_bits_entryid),
    .io_out_bits_awid(awreqArb_io_out_bits_awid),
    .io_out_bits_data(awreqArb_io_out_bits_data),
    .io_out_bits_mask(awreqArb_io_out_bits_mask),
    .io_out_bits_size(awreqArb_io_out_bits_size),
    .io_out_bits_len(awreqArb_io_out_bits_len)
  );
  Arbiter validreqArb ( // @[WriteStack.scala 62:27]
    .io_in_0_valid(validreqArb_io_in_0_valid),
    .io_in_0_bits_waddr(validreqArb_io_in_0_bits_waddr),
    .io_in_0_bits_entryid(validreqArb_io_in_0_bits_entryid),
    .io_in_0_bits_awid(validreqArb_io_in_0_bits_awid),
    .io_in_0_bits_data(validreqArb_io_in_0_bits_data),
    .io_in_0_bits_mask(validreqArb_io_in_0_bits_mask),
    .io_in_0_bits_size(validreqArb_io_in_0_bits_size),
    .io_in_0_bits_len(validreqArb_io_in_0_bits_len),
    .io_in_1_valid(validreqArb_io_in_1_valid),
    .io_in_1_bits_waddr(validreqArb_io_in_1_bits_waddr),
    .io_in_1_bits_entryid(validreqArb_io_in_1_bits_entryid),
    .io_in_1_bits_awid(validreqArb_io_in_1_bits_awid),
    .io_in_1_bits_data(validreqArb_io_in_1_bits_data),
    .io_in_1_bits_mask(validreqArb_io_in_1_bits_mask),
    .io_in_1_bits_size(validreqArb_io_in_1_bits_size),
    .io_in_1_bits_len(validreqArb_io_in_1_bits_len),
    .io_in_2_valid(validreqArb_io_in_2_valid),
    .io_in_2_bits_waddr(validreqArb_io_in_2_bits_waddr),
    .io_in_2_bits_entryid(validreqArb_io_in_2_bits_entryid),
    .io_in_2_bits_awid(validreqArb_io_in_2_bits_awid),
    .io_in_2_bits_data(validreqArb_io_in_2_bits_data),
    .io_in_2_bits_mask(validreqArb_io_in_2_bits_mask),
    .io_in_2_bits_size(validreqArb_io_in_2_bits_size),
    .io_in_2_bits_len(validreqArb_io_in_2_bits_len),
    .io_in_3_valid(validreqArb_io_in_3_valid),
    .io_in_3_bits_waddr(validreqArb_io_in_3_bits_waddr),
    .io_in_3_bits_entryid(validreqArb_io_in_3_bits_entryid),
    .io_in_3_bits_awid(validreqArb_io_in_3_bits_awid),
    .io_in_3_bits_data(validreqArb_io_in_3_bits_data),
    .io_in_3_bits_mask(validreqArb_io_in_3_bits_mask),
    .io_in_3_bits_size(validreqArb_io_in_3_bits_size),
    .io_in_3_bits_len(validreqArb_io_in_3_bits_len),
    .io_in_4_valid(validreqArb_io_in_4_valid),
    .io_in_4_bits_waddr(validreqArb_io_in_4_bits_waddr),
    .io_in_4_bits_entryid(validreqArb_io_in_4_bits_entryid),
    .io_in_4_bits_awid(validreqArb_io_in_4_bits_awid),
    .io_in_4_bits_data(validreqArb_io_in_4_bits_data),
    .io_in_4_bits_mask(validreqArb_io_in_4_bits_mask),
    .io_in_4_bits_size(validreqArb_io_in_4_bits_size),
    .io_in_4_bits_len(validreqArb_io_in_4_bits_len),
    .io_in_5_valid(validreqArb_io_in_5_valid),
    .io_in_5_bits_waddr(validreqArb_io_in_5_bits_waddr),
    .io_in_5_bits_entryid(validreqArb_io_in_5_bits_entryid),
    .io_in_5_bits_awid(validreqArb_io_in_5_bits_awid),
    .io_in_5_bits_data(validreqArb_io_in_5_bits_data),
    .io_in_5_bits_mask(validreqArb_io_in_5_bits_mask),
    .io_in_5_bits_size(validreqArb_io_in_5_bits_size),
    .io_in_5_bits_len(validreqArb_io_in_5_bits_len),
    .io_in_6_valid(validreqArb_io_in_6_valid),
    .io_in_6_bits_waddr(validreqArb_io_in_6_bits_waddr),
    .io_in_6_bits_entryid(validreqArb_io_in_6_bits_entryid),
    .io_in_6_bits_awid(validreqArb_io_in_6_bits_awid),
    .io_in_6_bits_data(validreqArb_io_in_6_bits_data),
    .io_in_6_bits_mask(validreqArb_io_in_6_bits_mask),
    .io_in_6_bits_size(validreqArb_io_in_6_bits_size),
    .io_in_6_bits_len(validreqArb_io_in_6_bits_len),
    .io_in_7_valid(validreqArb_io_in_7_valid),
    .io_in_7_bits_waddr(validreqArb_io_in_7_bits_waddr),
    .io_in_7_bits_entryid(validreqArb_io_in_7_bits_entryid),
    .io_in_7_bits_awid(validreqArb_io_in_7_bits_awid),
    .io_in_7_bits_data(validreqArb_io_in_7_bits_data),
    .io_in_7_bits_mask(validreqArb_io_in_7_bits_mask),
    .io_in_7_bits_size(validreqArb_io_in_7_bits_size),
    .io_in_7_bits_len(validreqArb_io_in_7_bits_len),
    .io_in_8_valid(validreqArb_io_in_8_valid),
    .io_in_8_bits_waddr(validreqArb_io_in_8_bits_waddr),
    .io_in_8_bits_entryid(validreqArb_io_in_8_bits_entryid),
    .io_in_8_bits_awid(validreqArb_io_in_8_bits_awid),
    .io_in_8_bits_data(validreqArb_io_in_8_bits_data),
    .io_in_8_bits_mask(validreqArb_io_in_8_bits_mask),
    .io_in_8_bits_size(validreqArb_io_in_8_bits_size),
    .io_in_8_bits_len(validreqArb_io_in_8_bits_len),
    .io_in_9_valid(validreqArb_io_in_9_valid),
    .io_in_9_bits_waddr(validreqArb_io_in_9_bits_waddr),
    .io_in_9_bits_entryid(validreqArb_io_in_9_bits_entryid),
    .io_in_9_bits_awid(validreqArb_io_in_9_bits_awid),
    .io_in_9_bits_data(validreqArb_io_in_9_bits_data),
    .io_in_9_bits_mask(validreqArb_io_in_9_bits_mask),
    .io_in_9_bits_size(validreqArb_io_in_9_bits_size),
    .io_in_9_bits_len(validreqArb_io_in_9_bits_len),
    .io_in_10_valid(validreqArb_io_in_10_valid),
    .io_in_10_bits_waddr(validreqArb_io_in_10_bits_waddr),
    .io_in_10_bits_entryid(validreqArb_io_in_10_bits_entryid),
    .io_in_10_bits_awid(validreqArb_io_in_10_bits_awid),
    .io_in_10_bits_data(validreqArb_io_in_10_bits_data),
    .io_in_10_bits_mask(validreqArb_io_in_10_bits_mask),
    .io_in_10_bits_size(validreqArb_io_in_10_bits_size),
    .io_in_10_bits_len(validreqArb_io_in_10_bits_len),
    .io_in_11_valid(validreqArb_io_in_11_valid),
    .io_in_11_bits_waddr(validreqArb_io_in_11_bits_waddr),
    .io_in_11_bits_entryid(validreqArb_io_in_11_bits_entryid),
    .io_in_11_bits_awid(validreqArb_io_in_11_bits_awid),
    .io_in_11_bits_data(validreqArb_io_in_11_bits_data),
    .io_in_11_bits_mask(validreqArb_io_in_11_bits_mask),
    .io_in_11_bits_size(validreqArb_io_in_11_bits_size),
    .io_in_11_bits_len(validreqArb_io_in_11_bits_len),
    .io_in_12_valid(validreqArb_io_in_12_valid),
    .io_in_12_bits_waddr(validreqArb_io_in_12_bits_waddr),
    .io_in_12_bits_entryid(validreqArb_io_in_12_bits_entryid),
    .io_in_12_bits_awid(validreqArb_io_in_12_bits_awid),
    .io_in_12_bits_data(validreqArb_io_in_12_bits_data),
    .io_in_12_bits_mask(validreqArb_io_in_12_bits_mask),
    .io_in_12_bits_size(validreqArb_io_in_12_bits_size),
    .io_in_12_bits_len(validreqArb_io_in_12_bits_len),
    .io_in_13_valid(validreqArb_io_in_13_valid),
    .io_in_13_bits_waddr(validreqArb_io_in_13_bits_waddr),
    .io_in_13_bits_entryid(validreqArb_io_in_13_bits_entryid),
    .io_in_13_bits_awid(validreqArb_io_in_13_bits_awid),
    .io_in_13_bits_data(validreqArb_io_in_13_bits_data),
    .io_in_13_bits_mask(validreqArb_io_in_13_bits_mask),
    .io_in_13_bits_size(validreqArb_io_in_13_bits_size),
    .io_in_13_bits_len(validreqArb_io_in_13_bits_len),
    .io_in_14_valid(validreqArb_io_in_14_valid),
    .io_in_14_bits_waddr(validreqArb_io_in_14_bits_waddr),
    .io_in_14_bits_entryid(validreqArb_io_in_14_bits_entryid),
    .io_in_14_bits_awid(validreqArb_io_in_14_bits_awid),
    .io_in_14_bits_data(validreqArb_io_in_14_bits_data),
    .io_in_14_bits_mask(validreqArb_io_in_14_bits_mask),
    .io_in_14_bits_size(validreqArb_io_in_14_bits_size),
    .io_in_14_bits_len(validreqArb_io_in_14_bits_len),
    .io_in_15_valid(validreqArb_io_in_15_valid),
    .io_in_15_bits_waddr(validreqArb_io_in_15_bits_waddr),
    .io_in_15_bits_entryid(validreqArb_io_in_15_bits_entryid),
    .io_in_15_bits_awid(validreqArb_io_in_15_bits_awid),
    .io_in_15_bits_data(validreqArb_io_in_15_bits_data),
    .io_in_15_bits_mask(validreqArb_io_in_15_bits_mask),
    .io_in_15_bits_size(validreqArb_io_in_15_bits_size),
    .io_in_15_bits_len(validreqArb_io_in_15_bits_len),
    .io_in_16_valid(validreqArb_io_in_16_valid),
    .io_in_16_bits_waddr(validreqArb_io_in_16_bits_waddr),
    .io_in_16_bits_entryid(validreqArb_io_in_16_bits_entryid),
    .io_in_16_bits_awid(validreqArb_io_in_16_bits_awid),
    .io_in_16_bits_data(validreqArb_io_in_16_bits_data),
    .io_in_16_bits_mask(validreqArb_io_in_16_bits_mask),
    .io_in_16_bits_size(validreqArb_io_in_16_bits_size),
    .io_in_16_bits_len(validreqArb_io_in_16_bits_len),
    .io_in_17_valid(validreqArb_io_in_17_valid),
    .io_in_17_bits_waddr(validreqArb_io_in_17_bits_waddr),
    .io_in_17_bits_entryid(validreqArb_io_in_17_bits_entryid),
    .io_in_17_bits_awid(validreqArb_io_in_17_bits_awid),
    .io_in_17_bits_data(validreqArb_io_in_17_bits_data),
    .io_in_17_bits_mask(validreqArb_io_in_17_bits_mask),
    .io_in_17_bits_size(validreqArb_io_in_17_bits_size),
    .io_in_17_bits_len(validreqArb_io_in_17_bits_len),
    .io_in_18_valid(validreqArb_io_in_18_valid),
    .io_in_18_bits_waddr(validreqArb_io_in_18_bits_waddr),
    .io_in_18_bits_entryid(validreqArb_io_in_18_bits_entryid),
    .io_in_18_bits_awid(validreqArb_io_in_18_bits_awid),
    .io_in_18_bits_data(validreqArb_io_in_18_bits_data),
    .io_in_18_bits_mask(validreqArb_io_in_18_bits_mask),
    .io_in_18_bits_size(validreqArb_io_in_18_bits_size),
    .io_in_18_bits_len(validreqArb_io_in_18_bits_len),
    .io_in_19_valid(validreqArb_io_in_19_valid),
    .io_in_19_bits_waddr(validreqArb_io_in_19_bits_waddr),
    .io_in_19_bits_entryid(validreqArb_io_in_19_bits_entryid),
    .io_in_19_bits_awid(validreqArb_io_in_19_bits_awid),
    .io_in_19_bits_data(validreqArb_io_in_19_bits_data),
    .io_in_19_bits_mask(validreqArb_io_in_19_bits_mask),
    .io_in_19_bits_size(validreqArb_io_in_19_bits_size),
    .io_in_19_bits_len(validreqArb_io_in_19_bits_len),
    .io_in_20_valid(validreqArb_io_in_20_valid),
    .io_in_20_bits_waddr(validreqArb_io_in_20_bits_waddr),
    .io_in_20_bits_entryid(validreqArb_io_in_20_bits_entryid),
    .io_in_20_bits_awid(validreqArb_io_in_20_bits_awid),
    .io_in_20_bits_data(validreqArb_io_in_20_bits_data),
    .io_in_20_bits_mask(validreqArb_io_in_20_bits_mask),
    .io_in_20_bits_size(validreqArb_io_in_20_bits_size),
    .io_in_20_bits_len(validreqArb_io_in_20_bits_len),
    .io_in_21_valid(validreqArb_io_in_21_valid),
    .io_in_21_bits_waddr(validreqArb_io_in_21_bits_waddr),
    .io_in_21_bits_entryid(validreqArb_io_in_21_bits_entryid),
    .io_in_21_bits_awid(validreqArb_io_in_21_bits_awid),
    .io_in_21_bits_data(validreqArb_io_in_21_bits_data),
    .io_in_21_bits_mask(validreqArb_io_in_21_bits_mask),
    .io_in_21_bits_size(validreqArb_io_in_21_bits_size),
    .io_in_21_bits_len(validreqArb_io_in_21_bits_len),
    .io_in_22_valid(validreqArb_io_in_22_valid),
    .io_in_22_bits_waddr(validreqArb_io_in_22_bits_waddr),
    .io_in_22_bits_entryid(validreqArb_io_in_22_bits_entryid),
    .io_in_22_bits_awid(validreqArb_io_in_22_bits_awid),
    .io_in_22_bits_data(validreqArb_io_in_22_bits_data),
    .io_in_22_bits_mask(validreqArb_io_in_22_bits_mask),
    .io_in_22_bits_size(validreqArb_io_in_22_bits_size),
    .io_in_22_bits_len(validreqArb_io_in_22_bits_len),
    .io_in_23_valid(validreqArb_io_in_23_valid),
    .io_in_23_bits_waddr(validreqArb_io_in_23_bits_waddr),
    .io_in_23_bits_entryid(validreqArb_io_in_23_bits_entryid),
    .io_in_23_bits_awid(validreqArb_io_in_23_bits_awid),
    .io_in_23_bits_data(validreqArb_io_in_23_bits_data),
    .io_in_23_bits_mask(validreqArb_io_in_23_bits_mask),
    .io_in_23_bits_size(validreqArb_io_in_23_bits_size),
    .io_in_23_bits_len(validreqArb_io_in_23_bits_len),
    .io_in_24_valid(validreqArb_io_in_24_valid),
    .io_in_24_bits_waddr(validreqArb_io_in_24_bits_waddr),
    .io_in_24_bits_entryid(validreqArb_io_in_24_bits_entryid),
    .io_in_24_bits_awid(validreqArb_io_in_24_bits_awid),
    .io_in_24_bits_data(validreqArb_io_in_24_bits_data),
    .io_in_24_bits_mask(validreqArb_io_in_24_bits_mask),
    .io_in_24_bits_size(validreqArb_io_in_24_bits_size),
    .io_in_24_bits_len(validreqArb_io_in_24_bits_len),
    .io_in_25_valid(validreqArb_io_in_25_valid),
    .io_in_25_bits_waddr(validreqArb_io_in_25_bits_waddr),
    .io_in_25_bits_entryid(validreqArb_io_in_25_bits_entryid),
    .io_in_25_bits_awid(validreqArb_io_in_25_bits_awid),
    .io_in_25_bits_data(validreqArb_io_in_25_bits_data),
    .io_in_25_bits_mask(validreqArb_io_in_25_bits_mask),
    .io_in_25_bits_size(validreqArb_io_in_25_bits_size),
    .io_in_25_bits_len(validreqArb_io_in_25_bits_len),
    .io_in_26_valid(validreqArb_io_in_26_valid),
    .io_in_26_bits_waddr(validreqArb_io_in_26_bits_waddr),
    .io_in_26_bits_entryid(validreqArb_io_in_26_bits_entryid),
    .io_in_26_bits_awid(validreqArb_io_in_26_bits_awid),
    .io_in_26_bits_data(validreqArb_io_in_26_bits_data),
    .io_in_26_bits_mask(validreqArb_io_in_26_bits_mask),
    .io_in_26_bits_size(validreqArb_io_in_26_bits_size),
    .io_in_26_bits_len(validreqArb_io_in_26_bits_len),
    .io_in_27_valid(validreqArb_io_in_27_valid),
    .io_in_27_bits_waddr(validreqArb_io_in_27_bits_waddr),
    .io_in_27_bits_entryid(validreqArb_io_in_27_bits_entryid),
    .io_in_27_bits_awid(validreqArb_io_in_27_bits_awid),
    .io_in_27_bits_data(validreqArb_io_in_27_bits_data),
    .io_in_27_bits_mask(validreqArb_io_in_27_bits_mask),
    .io_in_27_bits_size(validreqArb_io_in_27_bits_size),
    .io_in_27_bits_len(validreqArb_io_in_27_bits_len),
    .io_in_28_valid(validreqArb_io_in_28_valid),
    .io_in_28_bits_waddr(validreqArb_io_in_28_bits_waddr),
    .io_in_28_bits_entryid(validreqArb_io_in_28_bits_entryid),
    .io_in_28_bits_awid(validreqArb_io_in_28_bits_awid),
    .io_in_28_bits_data(validreqArb_io_in_28_bits_data),
    .io_in_28_bits_mask(validreqArb_io_in_28_bits_mask),
    .io_in_28_bits_size(validreqArb_io_in_28_bits_size),
    .io_in_28_bits_len(validreqArb_io_in_28_bits_len),
    .io_in_29_valid(validreqArb_io_in_29_valid),
    .io_in_29_bits_waddr(validreqArb_io_in_29_bits_waddr),
    .io_in_29_bits_entryid(validreqArb_io_in_29_bits_entryid),
    .io_in_29_bits_awid(validreqArb_io_in_29_bits_awid),
    .io_in_29_bits_data(validreqArb_io_in_29_bits_data),
    .io_in_29_bits_mask(validreqArb_io_in_29_bits_mask),
    .io_in_29_bits_size(validreqArb_io_in_29_bits_size),
    .io_in_29_bits_len(validreqArb_io_in_29_bits_len),
    .io_in_30_valid(validreqArb_io_in_30_valid),
    .io_in_30_bits_waddr(validreqArb_io_in_30_bits_waddr),
    .io_in_30_bits_entryid(validreqArb_io_in_30_bits_entryid),
    .io_in_30_bits_awid(validreqArb_io_in_30_bits_awid),
    .io_in_30_bits_data(validreqArb_io_in_30_bits_data),
    .io_in_30_bits_mask(validreqArb_io_in_30_bits_mask),
    .io_in_30_bits_size(validreqArb_io_in_30_bits_size),
    .io_in_30_bits_len(validreqArb_io_in_30_bits_len),
    .io_in_31_valid(validreqArb_io_in_31_valid),
    .io_in_31_bits_waddr(validreqArb_io_in_31_bits_waddr),
    .io_in_31_bits_entryid(validreqArb_io_in_31_bits_entryid),
    .io_in_31_bits_awid(validreqArb_io_in_31_bits_awid),
    .io_in_31_bits_data(validreqArb_io_in_31_bits_data),
    .io_in_31_bits_mask(validreqArb_io_in_31_bits_mask),
    .io_in_31_bits_size(validreqArb_io_in_31_bits_size),
    .io_in_31_bits_len(validreqArb_io_in_31_bits_len),
    .io_out_valid(validreqArb_io_out_valid),
    .io_out_bits_waddr(validreqArb_io_out_bits_waddr),
    .io_out_bits_entryid(validreqArb_io_out_bits_entryid),
    .io_out_bits_awid(validreqArb_io_out_bits_awid),
    .io_out_bits_data(validreqArb_io_out_bits_data),
    .io_out_bits_mask(validreqArb_io_out_bits_mask),
    .io_out_bits_size(validreqArb_io_out_bits_size),
    .io_out_bits_len(validreqArb_io_out_bits_len)
  );
  assign io_axiWriteReq_in_aw_ready = ~full; // @[WriteStack.scala 67:33]
  assign io_axiWriteReq_in_w_ready = |_canW_T_128; // @[WriteStack.scala 91:97]
  assign io_axiMenWriteReq_out_aw_valid = wreqArb_io_out_valid; // @[WriteStack.scala 181:34]
  assign io_axiMenWriteReq_out_aw_bits_id = wreqArb_io_out_bits_awid; // @[WriteStack.scala 182:36]
  assign io_axiMenWriteReq_out_aw_bits_addr = wreqArb_io_out_bits_waddr; // @[WriteStack.scala 183:38]
  assign io_axiMenWriteReq_out_aw_bits_len = wreqArb_io_out_bits_len; // @[WriteStack.scala 185:37]
  assign io_axiMenWriteReq_out_aw_bits_size = wreqArb_io_out_bits_size; // @[WriteStack.scala 184:38]
  assign io_axiMenWriteReq_out_aw_bits_burst = 2'h0; // @[WriteStack.scala 186:39]
  assign io_axiMenWriteReq_out_aw_bits_lock = 1'h0; // @[WriteStack.scala 187:38]
  assign io_axiMenWriteReq_out_aw_bits_cache = 4'h0; // @[WriteStack.scala 190:39]
  assign io_axiMenWriteReq_out_aw_bits_prot = 3'h0; // @[WriteStack.scala 188:38]
  assign io_axiMenWriteReq_out_aw_bits_qos = 4'h0; // @[WriteStack.scala 189:37]
  assign io_axiMenWriteReq_out_w_valid = awreqArb_io_out_valid; // @[WriteStack.scala 226:33]
  assign io_axiMenWriteReq_out_w_bits_data = awreqArb_io_out_bits_data; // @[WriteStack.scala 223:37]
  assign io_axiMenWriteReq_out_w_bits_strb = awreqArb_io_out_bits_mask; // @[WriteStack.scala 225:37]
  assign io_axiMenWriteReq_out_w_bits_last = 1'h1; // @[WriteStack.scala 224:37]
  assign io_axiMenWriteResp_in_b_ready = io_axiWriteResp_out_b_ready; // @[WriteStack.scala 252:33]
  assign io_axiWriteResp_out_b_valid = io_axiMenWriteResp_in_b_valid; // @[WriteStack.scala 251:31]
  assign io_axiWriteResp_out_b_bits_id = io_axiMenWriteResp_in_b_bits_id; // @[WriteStack.scala 253:30]
  assign io_axiWriteResp_out_b_bits_resp = io_axiMenWriteResp_in_b_bits_resp; // @[WriteStack.scala 253:30]
  assign io_validReq_in_valid = validreqArb_io_out_valid; // @[WriteStack.scala 136:24]
  assign io_validReq_in_bits_addr = validreqArb_io_out_bits_waddr; // @[WriteStack.scala 130:28]
  assign io_validReq_in_bits_source = {validreqArb_io_out_bits_entryid,validreqArb_io_out_bits_awid}; // @[Cat.scala 31:58]
  assign io_validResp_out_ready = |_canValid_T_64; // @[WriteStack.scala 162:88]
  assign wreqArb_io_in_0_valid = _canAW_T_3 & _canAW_T_4; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_0_bits_waddr = writeStack_0_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_entryid = writeStack_0_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_awid = writeStack_0_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_data = writeStack_0_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_mask = writeStack_0_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_size = writeStack_0_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_0_bits_len = writeStack_0_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_valid = _canAW_T_9 & _canAW_T_10; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_1_bits_waddr = writeStack_1_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_entryid = writeStack_1_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_awid = writeStack_1_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_data = writeStack_1_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_mask = writeStack_1_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_size = writeStack_1_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_1_bits_len = writeStack_1_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_valid = _canAW_T_15 & _canAW_T_16; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_2_bits_waddr = writeStack_2_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_entryid = writeStack_2_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_awid = writeStack_2_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_data = writeStack_2_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_mask = writeStack_2_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_size = writeStack_2_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_2_bits_len = writeStack_2_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_valid = _canAW_T_21 & _canAW_T_22; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_3_bits_waddr = writeStack_3_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_entryid = writeStack_3_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_awid = writeStack_3_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_data = writeStack_3_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_mask = writeStack_3_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_size = writeStack_3_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_3_bits_len = writeStack_3_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_valid = _canAW_T_27 & _canAW_T_28; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_4_bits_waddr = writeStack_4_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_entryid = writeStack_4_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_awid = writeStack_4_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_data = writeStack_4_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_mask = writeStack_4_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_size = writeStack_4_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_4_bits_len = writeStack_4_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_valid = _canAW_T_33 & _canAW_T_34; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_5_bits_waddr = writeStack_5_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_entryid = writeStack_5_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_awid = writeStack_5_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_data = writeStack_5_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_mask = writeStack_5_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_size = writeStack_5_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_5_bits_len = writeStack_5_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_valid = _canAW_T_39 & _canAW_T_40; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_6_bits_waddr = writeStack_6_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_entryid = writeStack_6_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_awid = writeStack_6_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_data = writeStack_6_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_mask = writeStack_6_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_size = writeStack_6_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_6_bits_len = writeStack_6_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_valid = _canAW_T_45 & _canAW_T_46; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_7_bits_waddr = writeStack_7_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_entryid = writeStack_7_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_awid = writeStack_7_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_data = writeStack_7_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_mask = writeStack_7_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_size = writeStack_7_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_7_bits_len = writeStack_7_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_valid = _canAW_T_51 & _canAW_T_52; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_8_bits_waddr = writeStack_8_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_entryid = writeStack_8_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_awid = writeStack_8_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_data = writeStack_8_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_mask = writeStack_8_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_size = writeStack_8_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_8_bits_len = writeStack_8_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_valid = _canAW_T_57 & _canAW_T_58; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_9_bits_waddr = writeStack_9_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_entryid = writeStack_9_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_awid = writeStack_9_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_data = writeStack_9_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_mask = writeStack_9_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_size = writeStack_9_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_9_bits_len = writeStack_9_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_valid = _canAW_T_63 & _canAW_T_64; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_10_bits_waddr = writeStack_10_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_entryid = writeStack_10_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_awid = writeStack_10_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_data = writeStack_10_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_mask = writeStack_10_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_size = writeStack_10_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_10_bits_len = writeStack_10_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_valid = _canAW_T_69 & _canAW_T_70; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_11_bits_waddr = writeStack_11_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_entryid = writeStack_11_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_awid = writeStack_11_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_data = writeStack_11_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_mask = writeStack_11_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_size = writeStack_11_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_11_bits_len = writeStack_11_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_valid = _canAW_T_75 & _canAW_T_76; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_12_bits_waddr = writeStack_12_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_entryid = writeStack_12_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_awid = writeStack_12_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_data = writeStack_12_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_mask = writeStack_12_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_size = writeStack_12_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_12_bits_len = writeStack_12_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_valid = _canAW_T_81 & _canAW_T_82; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_13_bits_waddr = writeStack_13_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_entryid = writeStack_13_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_awid = writeStack_13_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_data = writeStack_13_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_mask = writeStack_13_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_size = writeStack_13_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_13_bits_len = writeStack_13_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_valid = _canAW_T_87 & _canAW_T_88; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_14_bits_waddr = writeStack_14_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_entryid = writeStack_14_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_awid = writeStack_14_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_data = writeStack_14_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_mask = writeStack_14_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_size = writeStack_14_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_14_bits_len = writeStack_14_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_valid = _canAW_T_93 & _canAW_T_94; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_15_bits_waddr = writeStack_15_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_entryid = writeStack_15_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_awid = writeStack_15_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_data = writeStack_15_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_mask = writeStack_15_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_size = writeStack_15_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_15_bits_len = writeStack_15_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_valid = _canAW_T_99 & _canAW_T_100; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_16_bits_waddr = writeStack_16_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_entryid = writeStack_16_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_awid = writeStack_16_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_data = writeStack_16_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_mask = writeStack_16_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_size = writeStack_16_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_16_bits_len = writeStack_16_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_valid = _canAW_T_105 & _canAW_T_106; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_17_bits_waddr = writeStack_17_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_entryid = writeStack_17_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_awid = writeStack_17_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_data = writeStack_17_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_mask = writeStack_17_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_size = writeStack_17_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_17_bits_len = writeStack_17_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_valid = _canAW_T_111 & _canAW_T_112; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_18_bits_waddr = writeStack_18_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_entryid = writeStack_18_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_awid = writeStack_18_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_data = writeStack_18_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_mask = writeStack_18_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_size = writeStack_18_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_18_bits_len = writeStack_18_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_valid = _canAW_T_117 & _canAW_T_118; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_19_bits_waddr = writeStack_19_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_entryid = writeStack_19_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_awid = writeStack_19_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_data = writeStack_19_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_mask = writeStack_19_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_size = writeStack_19_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_19_bits_len = writeStack_19_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_valid = _canAW_T_123 & _canAW_T_124; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_20_bits_waddr = writeStack_20_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_entryid = writeStack_20_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_awid = writeStack_20_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_data = writeStack_20_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_mask = writeStack_20_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_size = writeStack_20_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_20_bits_len = writeStack_20_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_valid = _canAW_T_129 & _canAW_T_130; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_21_bits_waddr = writeStack_21_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_entryid = writeStack_21_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_awid = writeStack_21_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_data = writeStack_21_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_mask = writeStack_21_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_size = writeStack_21_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_21_bits_len = writeStack_21_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_valid = _canAW_T_135 & _canAW_T_136; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_22_bits_waddr = writeStack_22_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_entryid = writeStack_22_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_awid = writeStack_22_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_data = writeStack_22_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_mask = writeStack_22_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_size = writeStack_22_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_22_bits_len = writeStack_22_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_valid = _canAW_T_141 & _canAW_T_142; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_23_bits_waddr = writeStack_23_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_entryid = writeStack_23_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_awid = writeStack_23_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_data = writeStack_23_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_mask = writeStack_23_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_size = writeStack_23_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_23_bits_len = writeStack_23_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_valid = _canAW_T_147 & _canAW_T_148; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_24_bits_waddr = writeStack_24_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_entryid = writeStack_24_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_awid = writeStack_24_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_data = writeStack_24_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_mask = writeStack_24_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_size = writeStack_24_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_24_bits_len = writeStack_24_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_valid = _canAW_T_153 & _canAW_T_154; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_25_bits_waddr = writeStack_25_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_entryid = writeStack_25_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_awid = writeStack_25_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_data = writeStack_25_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_mask = writeStack_25_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_size = writeStack_25_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_25_bits_len = writeStack_25_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_valid = _canAW_T_159 & _canAW_T_160; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_26_bits_waddr = writeStack_26_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_entryid = writeStack_26_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_awid = writeStack_26_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_data = writeStack_26_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_mask = writeStack_26_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_size = writeStack_26_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_26_bits_len = writeStack_26_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_valid = _canAW_T_165 & _canAW_T_166; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_27_bits_waddr = writeStack_27_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_entryid = writeStack_27_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_awid = writeStack_27_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_data = writeStack_27_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_mask = writeStack_27_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_size = writeStack_27_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_27_bits_len = writeStack_27_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_valid = _canAW_T_171 & _canAW_T_172; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_28_bits_waddr = writeStack_28_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_entryid = writeStack_28_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_awid = writeStack_28_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_data = writeStack_28_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_mask = writeStack_28_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_size = writeStack_28_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_28_bits_len = writeStack_28_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_valid = _canAW_T_177 & _canAW_T_178; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_29_bits_waddr = writeStack_29_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_entryid = writeStack_29_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_awid = writeStack_29_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_data = writeStack_29_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_mask = writeStack_29_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_size = writeStack_29_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_29_bits_len = writeStack_29_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_valid = _canAW_T_183 & _canAW_T_184; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_30_bits_waddr = writeStack_30_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_entryid = writeStack_30_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_awid = writeStack_30_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_data = writeStack_30_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_mask = writeStack_30_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_size = writeStack_30_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_30_bits_len = writeStack_30_len; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_valid = _canAW_T_189 & _canAW_T_190; // @[WriteStack.scala 178:85]
  assign wreqArb_io_in_31_bits_waddr = writeStack_31_waddr; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_entryid = writeStack_31_entryid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_awid = writeStack_31_awid; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_data = writeStack_31_data; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_mask = writeStack_31_mask; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_size = writeStack_31_size; // @[WriteStack.scala 179:17]
  assign wreqArb_io_in_31_bits_len = writeStack_31_len; // @[WriteStack.scala 179:17]
  assign awreqArb_io_in_0_valid = _canMenW_T_3 & _canAW_T_4; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_0_bits_waddr = writeStack_0_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_entryid = writeStack_0_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_awid = writeStack_0_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_data = writeStack_0_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_mask = writeStack_0_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_size = writeStack_0_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_0_bits_len = writeStack_0_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_valid = _canMenW_T_9 & _canAW_T_10; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_1_bits_waddr = writeStack_1_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_entryid = writeStack_1_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_awid = writeStack_1_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_data = writeStack_1_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_mask = writeStack_1_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_size = writeStack_1_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_1_bits_len = writeStack_1_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_valid = _canMenW_T_15 & _canAW_T_16; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_2_bits_waddr = writeStack_2_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_entryid = writeStack_2_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_awid = writeStack_2_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_data = writeStack_2_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_mask = writeStack_2_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_size = writeStack_2_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_2_bits_len = writeStack_2_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_valid = _canMenW_T_21 & _canAW_T_22; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_3_bits_waddr = writeStack_3_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_entryid = writeStack_3_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_awid = writeStack_3_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_data = writeStack_3_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_mask = writeStack_3_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_size = writeStack_3_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_3_bits_len = writeStack_3_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_valid = _canMenW_T_27 & _canAW_T_28; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_4_bits_waddr = writeStack_4_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_entryid = writeStack_4_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_awid = writeStack_4_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_data = writeStack_4_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_mask = writeStack_4_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_size = writeStack_4_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_4_bits_len = writeStack_4_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_valid = _canMenW_T_33 & _canAW_T_34; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_5_bits_waddr = writeStack_5_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_entryid = writeStack_5_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_awid = writeStack_5_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_data = writeStack_5_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_mask = writeStack_5_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_size = writeStack_5_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_5_bits_len = writeStack_5_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_valid = _canMenW_T_39 & _canAW_T_40; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_6_bits_waddr = writeStack_6_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_entryid = writeStack_6_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_awid = writeStack_6_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_data = writeStack_6_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_mask = writeStack_6_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_size = writeStack_6_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_6_bits_len = writeStack_6_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_valid = _canMenW_T_45 & _canAW_T_46; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_7_bits_waddr = writeStack_7_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_entryid = writeStack_7_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_awid = writeStack_7_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_data = writeStack_7_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_mask = writeStack_7_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_size = writeStack_7_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_7_bits_len = writeStack_7_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_valid = _canMenW_T_51 & _canAW_T_52; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_8_bits_waddr = writeStack_8_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_entryid = writeStack_8_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_awid = writeStack_8_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_data = writeStack_8_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_mask = writeStack_8_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_size = writeStack_8_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_8_bits_len = writeStack_8_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_valid = _canMenW_T_57 & _canAW_T_58; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_9_bits_waddr = writeStack_9_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_entryid = writeStack_9_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_awid = writeStack_9_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_data = writeStack_9_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_mask = writeStack_9_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_size = writeStack_9_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_9_bits_len = writeStack_9_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_valid = _canMenW_T_63 & _canAW_T_64; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_10_bits_waddr = writeStack_10_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_entryid = writeStack_10_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_awid = writeStack_10_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_data = writeStack_10_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_mask = writeStack_10_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_size = writeStack_10_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_10_bits_len = writeStack_10_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_valid = _canMenW_T_69 & _canAW_T_70; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_11_bits_waddr = writeStack_11_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_entryid = writeStack_11_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_awid = writeStack_11_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_data = writeStack_11_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_mask = writeStack_11_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_size = writeStack_11_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_11_bits_len = writeStack_11_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_valid = _canMenW_T_75 & _canAW_T_76; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_12_bits_waddr = writeStack_12_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_entryid = writeStack_12_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_awid = writeStack_12_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_data = writeStack_12_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_mask = writeStack_12_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_size = writeStack_12_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_12_bits_len = writeStack_12_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_valid = _canMenW_T_81 & _canAW_T_82; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_13_bits_waddr = writeStack_13_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_entryid = writeStack_13_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_awid = writeStack_13_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_data = writeStack_13_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_mask = writeStack_13_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_size = writeStack_13_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_13_bits_len = writeStack_13_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_valid = _canMenW_T_87 & _canAW_T_88; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_14_bits_waddr = writeStack_14_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_entryid = writeStack_14_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_awid = writeStack_14_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_data = writeStack_14_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_mask = writeStack_14_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_size = writeStack_14_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_14_bits_len = writeStack_14_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_valid = _canMenW_T_93 & _canAW_T_94; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_15_bits_waddr = writeStack_15_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_entryid = writeStack_15_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_awid = writeStack_15_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_data = writeStack_15_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_mask = writeStack_15_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_size = writeStack_15_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_15_bits_len = writeStack_15_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_valid = _canMenW_T_99 & _canAW_T_100; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_16_bits_waddr = writeStack_16_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_entryid = writeStack_16_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_awid = writeStack_16_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_data = writeStack_16_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_mask = writeStack_16_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_size = writeStack_16_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_16_bits_len = writeStack_16_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_valid = _canMenW_T_105 & _canAW_T_106; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_17_bits_waddr = writeStack_17_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_entryid = writeStack_17_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_awid = writeStack_17_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_data = writeStack_17_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_mask = writeStack_17_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_size = writeStack_17_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_17_bits_len = writeStack_17_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_valid = _canMenW_T_111 & _canAW_T_112; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_18_bits_waddr = writeStack_18_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_entryid = writeStack_18_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_awid = writeStack_18_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_data = writeStack_18_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_mask = writeStack_18_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_size = writeStack_18_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_18_bits_len = writeStack_18_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_valid = _canMenW_T_117 & _canAW_T_118; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_19_bits_waddr = writeStack_19_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_entryid = writeStack_19_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_awid = writeStack_19_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_data = writeStack_19_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_mask = writeStack_19_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_size = writeStack_19_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_19_bits_len = writeStack_19_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_valid = _canMenW_T_123 & _canAW_T_124; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_20_bits_waddr = writeStack_20_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_entryid = writeStack_20_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_awid = writeStack_20_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_data = writeStack_20_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_mask = writeStack_20_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_size = writeStack_20_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_20_bits_len = writeStack_20_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_valid = _canMenW_T_129 & _canAW_T_130; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_21_bits_waddr = writeStack_21_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_entryid = writeStack_21_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_awid = writeStack_21_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_data = writeStack_21_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_mask = writeStack_21_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_size = writeStack_21_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_21_bits_len = writeStack_21_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_valid = _canMenW_T_135 & _canAW_T_136; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_22_bits_waddr = writeStack_22_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_entryid = writeStack_22_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_awid = writeStack_22_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_data = writeStack_22_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_mask = writeStack_22_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_size = writeStack_22_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_22_bits_len = writeStack_22_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_valid = _canMenW_T_141 & _canAW_T_142; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_23_bits_waddr = writeStack_23_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_entryid = writeStack_23_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_awid = writeStack_23_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_data = writeStack_23_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_mask = writeStack_23_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_size = writeStack_23_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_23_bits_len = writeStack_23_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_valid = _canMenW_T_147 & _canAW_T_148; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_24_bits_waddr = writeStack_24_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_entryid = writeStack_24_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_awid = writeStack_24_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_data = writeStack_24_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_mask = writeStack_24_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_size = writeStack_24_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_24_bits_len = writeStack_24_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_valid = _canMenW_T_153 & _canAW_T_154; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_25_bits_waddr = writeStack_25_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_entryid = writeStack_25_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_awid = writeStack_25_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_data = writeStack_25_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_mask = writeStack_25_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_size = writeStack_25_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_25_bits_len = writeStack_25_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_valid = _canMenW_T_159 & _canAW_T_160; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_26_bits_waddr = writeStack_26_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_entryid = writeStack_26_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_awid = writeStack_26_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_data = writeStack_26_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_mask = writeStack_26_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_size = writeStack_26_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_26_bits_len = writeStack_26_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_valid = _canMenW_T_165 & _canAW_T_166; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_27_bits_waddr = writeStack_27_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_entryid = writeStack_27_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_awid = writeStack_27_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_data = writeStack_27_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_mask = writeStack_27_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_size = writeStack_27_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_27_bits_len = writeStack_27_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_valid = _canMenW_T_171 & _canAW_T_172; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_28_bits_waddr = writeStack_28_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_entryid = writeStack_28_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_awid = writeStack_28_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_data = writeStack_28_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_mask = writeStack_28_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_size = writeStack_28_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_28_bits_len = writeStack_28_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_valid = _canMenW_T_177 & _canAW_T_178; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_29_bits_waddr = writeStack_29_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_entryid = writeStack_29_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_awid = writeStack_29_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_data = writeStack_29_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_mask = writeStack_29_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_size = writeStack_29_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_29_bits_len = writeStack_29_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_valid = _canMenW_T_183 & _canAW_T_184; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_30_bits_waddr = writeStack_30_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_entryid = writeStack_30_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_awid = writeStack_30_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_data = writeStack_30_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_mask = writeStack_30_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_size = writeStack_30_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_30_bits_len = writeStack_30_len; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_valid = _canMenW_T_189 & _canAW_T_190; // @[WriteStack.scala 220:85]
  assign awreqArb_io_in_31_bits_waddr = writeStack_31_waddr; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_entryid = writeStack_31_entryid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_awid = writeStack_31_awid; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_data = writeStack_31_data; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_mask = writeStack_31_mask; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_size = writeStack_31_size; // @[WriteStack.scala 221:17]
  assign awreqArb_io_in_31_bits_len = writeStack_31_len; // @[WriteStack.scala 221:17]
  assign validreqArb_io_in_0_valid = _hasValid_T_2 & writeStack_0_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_0_bits_waddr = writeStack_0_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_entryid = writeStack_0_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_awid = writeStack_0_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_data = writeStack_0_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_mask = writeStack_0_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_size = writeStack_0_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_0_bits_len = writeStack_0_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_valid = _hasValid_T_5 & writeStack_1_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_1_bits_waddr = writeStack_1_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_entryid = writeStack_1_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_awid = writeStack_1_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_data = writeStack_1_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_mask = writeStack_1_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_size = writeStack_1_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_1_bits_len = writeStack_1_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_valid = _hasValid_T_8 & writeStack_2_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_2_bits_waddr = writeStack_2_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_entryid = writeStack_2_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_awid = writeStack_2_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_data = writeStack_2_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_mask = writeStack_2_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_size = writeStack_2_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_2_bits_len = writeStack_2_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_valid = _hasValid_T_11 & writeStack_3_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_3_bits_waddr = writeStack_3_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_entryid = writeStack_3_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_awid = writeStack_3_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_data = writeStack_3_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_mask = writeStack_3_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_size = writeStack_3_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_3_bits_len = writeStack_3_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_valid = _hasValid_T_14 & writeStack_4_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_4_bits_waddr = writeStack_4_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_entryid = writeStack_4_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_awid = writeStack_4_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_data = writeStack_4_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_mask = writeStack_4_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_size = writeStack_4_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_4_bits_len = writeStack_4_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_valid = _hasValid_T_17 & writeStack_5_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_5_bits_waddr = writeStack_5_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_entryid = writeStack_5_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_awid = writeStack_5_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_data = writeStack_5_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_mask = writeStack_5_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_size = writeStack_5_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_5_bits_len = writeStack_5_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_valid = _hasValid_T_20 & writeStack_6_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_6_bits_waddr = writeStack_6_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_entryid = writeStack_6_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_awid = writeStack_6_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_data = writeStack_6_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_mask = writeStack_6_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_size = writeStack_6_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_6_bits_len = writeStack_6_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_valid = _hasValid_T_23 & writeStack_7_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_7_bits_waddr = writeStack_7_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_entryid = writeStack_7_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_awid = writeStack_7_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_data = writeStack_7_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_mask = writeStack_7_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_size = writeStack_7_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_7_bits_len = writeStack_7_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_valid = _hasValid_T_26 & writeStack_8_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_8_bits_waddr = writeStack_8_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_entryid = writeStack_8_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_awid = writeStack_8_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_data = writeStack_8_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_mask = writeStack_8_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_size = writeStack_8_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_8_bits_len = writeStack_8_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_valid = _hasValid_T_29 & writeStack_9_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_9_bits_waddr = writeStack_9_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_entryid = writeStack_9_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_awid = writeStack_9_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_data = writeStack_9_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_mask = writeStack_9_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_size = writeStack_9_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_9_bits_len = writeStack_9_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_valid = _hasValid_T_32 & writeStack_10_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_10_bits_waddr = writeStack_10_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_entryid = writeStack_10_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_awid = writeStack_10_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_data = writeStack_10_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_mask = writeStack_10_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_size = writeStack_10_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_10_bits_len = writeStack_10_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_valid = _hasValid_T_35 & writeStack_11_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_11_bits_waddr = writeStack_11_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_entryid = writeStack_11_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_awid = writeStack_11_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_data = writeStack_11_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_mask = writeStack_11_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_size = writeStack_11_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_11_bits_len = writeStack_11_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_valid = _hasValid_T_38 & writeStack_12_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_12_bits_waddr = writeStack_12_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_entryid = writeStack_12_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_awid = writeStack_12_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_data = writeStack_12_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_mask = writeStack_12_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_size = writeStack_12_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_12_bits_len = writeStack_12_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_valid = _hasValid_T_41 & writeStack_13_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_13_bits_waddr = writeStack_13_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_entryid = writeStack_13_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_awid = writeStack_13_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_data = writeStack_13_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_mask = writeStack_13_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_size = writeStack_13_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_13_bits_len = writeStack_13_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_valid = _hasValid_T_44 & writeStack_14_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_14_bits_waddr = writeStack_14_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_entryid = writeStack_14_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_awid = writeStack_14_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_data = writeStack_14_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_mask = writeStack_14_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_size = writeStack_14_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_14_bits_len = writeStack_14_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_valid = _hasValid_T_47 & writeStack_15_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_15_bits_waddr = writeStack_15_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_entryid = writeStack_15_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_awid = writeStack_15_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_data = writeStack_15_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_mask = writeStack_15_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_size = writeStack_15_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_15_bits_len = writeStack_15_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_valid = _hasValid_T_50 & writeStack_16_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_16_bits_waddr = writeStack_16_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_entryid = writeStack_16_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_awid = writeStack_16_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_data = writeStack_16_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_mask = writeStack_16_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_size = writeStack_16_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_16_bits_len = writeStack_16_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_valid = _hasValid_T_53 & writeStack_17_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_17_bits_waddr = writeStack_17_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_entryid = writeStack_17_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_awid = writeStack_17_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_data = writeStack_17_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_mask = writeStack_17_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_size = writeStack_17_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_17_bits_len = writeStack_17_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_valid = _hasValid_T_56 & writeStack_18_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_18_bits_waddr = writeStack_18_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_entryid = writeStack_18_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_awid = writeStack_18_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_data = writeStack_18_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_mask = writeStack_18_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_size = writeStack_18_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_18_bits_len = writeStack_18_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_valid = _hasValid_T_59 & writeStack_19_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_19_bits_waddr = writeStack_19_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_entryid = writeStack_19_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_awid = writeStack_19_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_data = writeStack_19_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_mask = writeStack_19_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_size = writeStack_19_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_19_bits_len = writeStack_19_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_valid = _hasValid_T_62 & writeStack_20_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_20_bits_waddr = writeStack_20_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_entryid = writeStack_20_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_awid = writeStack_20_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_data = writeStack_20_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_mask = writeStack_20_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_size = writeStack_20_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_20_bits_len = writeStack_20_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_valid = _hasValid_T_65 & writeStack_21_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_21_bits_waddr = writeStack_21_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_entryid = writeStack_21_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_awid = writeStack_21_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_data = writeStack_21_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_mask = writeStack_21_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_size = writeStack_21_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_21_bits_len = writeStack_21_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_valid = _hasValid_T_68 & writeStack_22_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_22_bits_waddr = writeStack_22_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_entryid = writeStack_22_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_awid = writeStack_22_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_data = writeStack_22_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_mask = writeStack_22_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_size = writeStack_22_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_22_bits_len = writeStack_22_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_valid = _hasValid_T_71 & writeStack_23_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_23_bits_waddr = writeStack_23_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_entryid = writeStack_23_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_awid = writeStack_23_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_data = writeStack_23_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_mask = writeStack_23_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_size = writeStack_23_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_23_bits_len = writeStack_23_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_valid = _hasValid_T_74 & writeStack_24_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_24_bits_waddr = writeStack_24_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_entryid = writeStack_24_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_awid = writeStack_24_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_data = writeStack_24_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_mask = writeStack_24_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_size = writeStack_24_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_24_bits_len = writeStack_24_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_valid = _hasValid_T_77 & writeStack_25_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_25_bits_waddr = writeStack_25_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_entryid = writeStack_25_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_awid = writeStack_25_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_data = writeStack_25_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_mask = writeStack_25_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_size = writeStack_25_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_25_bits_len = writeStack_25_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_valid = _hasValid_T_80 & writeStack_26_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_26_bits_waddr = writeStack_26_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_entryid = writeStack_26_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_awid = writeStack_26_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_data = writeStack_26_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_mask = writeStack_26_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_size = writeStack_26_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_26_bits_len = writeStack_26_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_valid = _hasValid_T_83 & writeStack_27_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_27_bits_waddr = writeStack_27_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_entryid = writeStack_27_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_awid = writeStack_27_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_data = writeStack_27_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_mask = writeStack_27_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_size = writeStack_27_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_27_bits_len = writeStack_27_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_valid = _hasValid_T_86 & writeStack_28_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_28_bits_waddr = writeStack_28_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_entryid = writeStack_28_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_awid = writeStack_28_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_data = writeStack_28_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_mask = writeStack_28_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_size = writeStack_28_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_28_bits_len = writeStack_28_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_valid = _hasValid_T_89 & writeStack_29_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_29_bits_waddr = writeStack_29_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_entryid = writeStack_29_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_awid = writeStack_29_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_data = writeStack_29_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_mask = writeStack_29_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_size = writeStack_29_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_29_bits_len = writeStack_29_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_valid = _hasValid_T_92 & writeStack_30_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_30_bits_waddr = writeStack_30_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_entryid = writeStack_30_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_awid = writeStack_30_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_data = writeStack_30_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_mask = writeStack_30_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_size = writeStack_30_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_30_bits_len = writeStack_30_len; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_valid = _hasValid_T_95 & writeStack_31_wvalid; // @[WriteStack.scala 126:74]
  assign validreqArb_io_in_31_bits_waddr = writeStack_31_waddr; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_entryid = writeStack_31_entryid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_awid = writeStack_31_awid; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_data = writeStack_31_data; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_mask = writeStack_31_mask; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_size = writeStack_31_size; // @[WriteStack.scala 127:17]
  assign validreqArb_io_in_31_bits_len = writeStack_31_len; // @[WriteStack.scala 127:17]
  always @(posedge clock) begin
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_5) begin // @[WriteStack.scala 233:15]
        writeStack_0_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_0_wvalid <= _GEN_288;
      end
    end else begin
      writeStack_0_wvalid <= _GEN_288;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h0 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_0_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_0_wstatus <= _GEN_2432[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h0 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_0_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_0_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h0 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_0_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_5) begin // @[WriteStack.scala 233:15]
        writeStack_0_entryFifoid <= _writeStack_0_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_609) begin // @[WriteStack.scala 240:15]
        writeStack_0_entryFifoid <= _writeStack_0_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_0_entryFifoid <= _GEN_1440;
      end
    end else begin
      writeStack_0_entryFifoid <= _GEN_1440;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_1 & _hasValid_T_1) begin // @[WriteStack.scala 151:84]
        writeStack_0_validFifoId <= _writeStack_0_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_1) begin // @[WriteStack.scala 154:65]
        writeStack_0_validFifoId <= _writeStack_0_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_0_validFifoId <= _GEN_1088;
      end
    end else begin
      writeStack_0_validFifoId <= _GEN_1088;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_3) begin // @[WriteStack.scala 109:76]
        writeStack_0_waitWFifoId <= _writeStack_0_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_1) begin // @[WriteStack.scala 115:15]
        writeStack_0_waitWFifoId <= _writeStack_0_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_0_waitWFifoId <= _GEN_672;
      end
    end else begin
      writeStack_0_waitWFifoId <= _GEN_672;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_3) begin // @[WriteStack.scala 109:76]
        writeStack_0_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_3) begin // @[WriteStack.scala 109:76]
        writeStack_0_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_0_validStatus <= _GEN_2433[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h0 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_0_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_0_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h0 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_0_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_11) begin // @[WriteStack.scala 233:15]
        writeStack_1_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_1_wvalid <= _GEN_289;
      end
    end else begin
      writeStack_1_wvalid <= _GEN_289;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_1_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_1_wstatus <= _GEN_2434[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_1_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_1_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_1_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_11) begin // @[WriteStack.scala 233:15]
        writeStack_1_entryFifoid <= _writeStack_1_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_617) begin // @[WriteStack.scala 240:15]
        writeStack_1_entryFifoid <= _writeStack_1_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_1_entryFifoid <= _GEN_1441;
      end
    end else begin
      writeStack_1_entryFifoid <= _GEN_1441;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_3 & _hasValid_T_4) begin // @[WriteStack.scala 151:84]
        writeStack_1_validFifoId <= _writeStack_1_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_3) begin // @[WriteStack.scala 154:65]
        writeStack_1_validFifoId <= _writeStack_1_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_1_validFifoId <= _GEN_1089;
      end
    end else begin
      writeStack_1_validFifoId <= _GEN_1089;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_7) begin // @[WriteStack.scala 109:76]
        writeStack_1_waitWFifoId <= _writeStack_1_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_5) begin // @[WriteStack.scala 115:15]
        writeStack_1_waitWFifoId <= _writeStack_1_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_1_waitWFifoId <= _GEN_673;
      end
    end else begin
      writeStack_1_waitWFifoId <= _GEN_673;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_7) begin // @[WriteStack.scala 109:76]
        writeStack_1_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_7) begin // @[WriteStack.scala 109:76]
        writeStack_1_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_1_validStatus <= _GEN_2435[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_1_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_1_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_1_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_17) begin // @[WriteStack.scala 233:15]
        writeStack_2_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_2_wvalid <= _GEN_290;
      end
    end else begin
      writeStack_2_wvalid <= _GEN_290;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h2 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_2_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_2_wstatus <= _GEN_2436[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h2 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_2_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_2_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h2 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_2_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_17) begin // @[WriteStack.scala 233:15]
        writeStack_2_entryFifoid <= _writeStack_2_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_625) begin // @[WriteStack.scala 240:15]
        writeStack_2_entryFifoid <= _writeStack_2_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_2_entryFifoid <= _GEN_1442;
      end
    end else begin
      writeStack_2_entryFifoid <= _GEN_1442;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_5 & _hasValid_T_7) begin // @[WriteStack.scala 151:84]
        writeStack_2_validFifoId <= _writeStack_2_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_5) begin // @[WriteStack.scala 154:65]
        writeStack_2_validFifoId <= _writeStack_2_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_2_validFifoId <= _GEN_1090;
      end
    end else begin
      writeStack_2_validFifoId <= _GEN_1090;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_11) begin // @[WriteStack.scala 109:76]
        writeStack_2_waitWFifoId <= _writeStack_2_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_9) begin // @[WriteStack.scala 115:15]
        writeStack_2_waitWFifoId <= _writeStack_2_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_2_waitWFifoId <= _GEN_674;
      end
    end else begin
      writeStack_2_waitWFifoId <= _GEN_674;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_11) begin // @[WriteStack.scala 109:76]
        writeStack_2_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_11) begin // @[WriteStack.scala 109:76]
        writeStack_2_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_2_validStatus <= _GEN_2437[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h2 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_2_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_2_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h2 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_2_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_23) begin // @[WriteStack.scala 233:15]
        writeStack_3_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_3_wvalid <= _GEN_291;
      end
    end else begin
      writeStack_3_wvalid <= _GEN_291;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h3 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_3_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_3_wstatus <= _GEN_2438[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h3 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_3_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_3_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h3 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_3_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_23) begin // @[WriteStack.scala 233:15]
        writeStack_3_entryFifoid <= _writeStack_3_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_633) begin // @[WriteStack.scala 240:15]
        writeStack_3_entryFifoid <= _writeStack_3_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_3_entryFifoid <= _GEN_1443;
      end
    end else begin
      writeStack_3_entryFifoid <= _GEN_1443;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_7 & _hasValid_T_10) begin // @[WriteStack.scala 151:84]
        writeStack_3_validFifoId <= _writeStack_3_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_7) begin // @[WriteStack.scala 154:65]
        writeStack_3_validFifoId <= _writeStack_3_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_3_validFifoId <= _GEN_1091;
      end
    end else begin
      writeStack_3_validFifoId <= _GEN_1091;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_15) begin // @[WriteStack.scala 109:76]
        writeStack_3_waitWFifoId <= _writeStack_3_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_13) begin // @[WriteStack.scala 115:15]
        writeStack_3_waitWFifoId <= _writeStack_3_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_3_waitWFifoId <= _GEN_675;
      end
    end else begin
      writeStack_3_waitWFifoId <= _GEN_675;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_15) begin // @[WriteStack.scala 109:76]
        writeStack_3_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_15) begin // @[WriteStack.scala 109:76]
        writeStack_3_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_3_validStatus <= _GEN_2439[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h3 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_3_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_3_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h3 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_3_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_29) begin // @[WriteStack.scala 233:15]
        writeStack_4_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_4_wvalid <= _GEN_292;
      end
    end else begin
      writeStack_4_wvalid <= _GEN_292;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h4 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_4_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_4_wstatus <= _GEN_2440[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h4 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_4_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_4_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h4 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_4_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_29) begin // @[WriteStack.scala 233:15]
        writeStack_4_entryFifoid <= _writeStack_4_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_641) begin // @[WriteStack.scala 240:15]
        writeStack_4_entryFifoid <= _writeStack_4_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_4_entryFifoid <= _GEN_1444;
      end
    end else begin
      writeStack_4_entryFifoid <= _GEN_1444;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_9 & _hasValid_T_13) begin // @[WriteStack.scala 151:84]
        writeStack_4_validFifoId <= _writeStack_4_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_9) begin // @[WriteStack.scala 154:65]
        writeStack_4_validFifoId <= _writeStack_4_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_4_validFifoId <= _GEN_1092;
      end
    end else begin
      writeStack_4_validFifoId <= _GEN_1092;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_19) begin // @[WriteStack.scala 109:76]
        writeStack_4_waitWFifoId <= _writeStack_4_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_17) begin // @[WriteStack.scala 115:15]
        writeStack_4_waitWFifoId <= _writeStack_4_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_4_waitWFifoId <= _GEN_676;
      end
    end else begin
      writeStack_4_waitWFifoId <= _GEN_676;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_19) begin // @[WriteStack.scala 109:76]
        writeStack_4_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_19) begin // @[WriteStack.scala 109:76]
        writeStack_4_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_4_validStatus <= _GEN_2441[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h4 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_4_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_4_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h4 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_4_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_35) begin // @[WriteStack.scala 233:15]
        writeStack_5_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_5_wvalid <= _GEN_293;
      end
    end else begin
      writeStack_5_wvalid <= _GEN_293;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h5 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_5_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_5_wstatus <= _GEN_2442[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h5 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_5_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_5_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h5 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_5_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_35) begin // @[WriteStack.scala 233:15]
        writeStack_5_entryFifoid <= _writeStack_5_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_649) begin // @[WriteStack.scala 240:15]
        writeStack_5_entryFifoid <= _writeStack_5_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_5_entryFifoid <= _GEN_1445;
      end
    end else begin
      writeStack_5_entryFifoid <= _GEN_1445;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_11 & _hasValid_T_16) begin // @[WriteStack.scala 151:84]
        writeStack_5_validFifoId <= _writeStack_5_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_11) begin // @[WriteStack.scala 154:65]
        writeStack_5_validFifoId <= _writeStack_5_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_5_validFifoId <= _GEN_1093;
      end
    end else begin
      writeStack_5_validFifoId <= _GEN_1093;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_23) begin // @[WriteStack.scala 109:76]
        writeStack_5_waitWFifoId <= _writeStack_5_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_21) begin // @[WriteStack.scala 115:15]
        writeStack_5_waitWFifoId <= _writeStack_5_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_5_waitWFifoId <= _GEN_677;
      end
    end else begin
      writeStack_5_waitWFifoId <= _GEN_677;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_23) begin // @[WriteStack.scala 109:76]
        writeStack_5_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_23) begin // @[WriteStack.scala 109:76]
        writeStack_5_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_5_validStatus <= _GEN_2443[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h5 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_5_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_5_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h5 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_5_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_41) begin // @[WriteStack.scala 233:15]
        writeStack_6_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_6_wvalid <= _GEN_294;
      end
    end else begin
      writeStack_6_wvalid <= _GEN_294;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h6 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_6_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_6_wstatus <= _GEN_2444[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h6 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_6_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_6_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h6 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_6_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_41) begin // @[WriteStack.scala 233:15]
        writeStack_6_entryFifoid <= _writeStack_6_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_657) begin // @[WriteStack.scala 240:15]
        writeStack_6_entryFifoid <= _writeStack_6_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_6_entryFifoid <= _GEN_1446;
      end
    end else begin
      writeStack_6_entryFifoid <= _GEN_1446;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_13 & _hasValid_T_19) begin // @[WriteStack.scala 151:84]
        writeStack_6_validFifoId <= _writeStack_6_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_13) begin // @[WriteStack.scala 154:65]
        writeStack_6_validFifoId <= _writeStack_6_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_6_validFifoId <= _GEN_1094;
      end
    end else begin
      writeStack_6_validFifoId <= _GEN_1094;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_27) begin // @[WriteStack.scala 109:76]
        writeStack_6_waitWFifoId <= _writeStack_6_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_25) begin // @[WriteStack.scala 115:15]
        writeStack_6_waitWFifoId <= _writeStack_6_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_6_waitWFifoId <= _GEN_678;
      end
    end else begin
      writeStack_6_waitWFifoId <= _GEN_678;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_27) begin // @[WriteStack.scala 109:76]
        writeStack_6_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_27) begin // @[WriteStack.scala 109:76]
        writeStack_6_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_6_validStatus <= _GEN_2445[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h6 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_6_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_6_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h6 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_6_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_47) begin // @[WriteStack.scala 233:15]
        writeStack_7_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_7_wvalid <= _GEN_295;
      end
    end else begin
      writeStack_7_wvalid <= _GEN_295;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h7 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_7_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_7_wstatus <= _GEN_2446[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h7 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_7_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_7_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h7 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_7_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_47) begin // @[WriteStack.scala 233:15]
        writeStack_7_entryFifoid <= _writeStack_7_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_665) begin // @[WriteStack.scala 240:15]
        writeStack_7_entryFifoid <= _writeStack_7_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_7_entryFifoid <= _GEN_1447;
      end
    end else begin
      writeStack_7_entryFifoid <= _GEN_1447;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_15 & _hasValid_T_22) begin // @[WriteStack.scala 151:84]
        writeStack_7_validFifoId <= _writeStack_7_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_15) begin // @[WriteStack.scala 154:65]
        writeStack_7_validFifoId <= _writeStack_7_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_7_validFifoId <= _GEN_1095;
      end
    end else begin
      writeStack_7_validFifoId <= _GEN_1095;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_31) begin // @[WriteStack.scala 109:76]
        writeStack_7_waitWFifoId <= _writeStack_7_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_29) begin // @[WriteStack.scala 115:15]
        writeStack_7_waitWFifoId <= _writeStack_7_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_7_waitWFifoId <= _GEN_679;
      end
    end else begin
      writeStack_7_waitWFifoId <= _GEN_679;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_31) begin // @[WriteStack.scala 109:76]
        writeStack_7_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_31) begin // @[WriteStack.scala 109:76]
        writeStack_7_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_7_validStatus <= _GEN_2447[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h7 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_7_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_7_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h7 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_7_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_53) begin // @[WriteStack.scala 233:15]
        writeStack_8_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_8_wvalid <= _GEN_296;
      end
    end else begin
      writeStack_8_wvalid <= _GEN_296;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h8 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_8_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_8_wstatus <= _GEN_2448[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h8 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_8_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_8_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h8 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_8_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_53) begin // @[WriteStack.scala 233:15]
        writeStack_8_entryFifoid <= _writeStack_8_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_673) begin // @[WriteStack.scala 240:15]
        writeStack_8_entryFifoid <= _writeStack_8_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_8_entryFifoid <= _GEN_1448;
      end
    end else begin
      writeStack_8_entryFifoid <= _GEN_1448;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_17 & _hasValid_T_25) begin // @[WriteStack.scala 151:84]
        writeStack_8_validFifoId <= _writeStack_8_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_17) begin // @[WriteStack.scala 154:65]
        writeStack_8_validFifoId <= _writeStack_8_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_8_validFifoId <= _GEN_1096;
      end
    end else begin
      writeStack_8_validFifoId <= _GEN_1096;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_35) begin // @[WriteStack.scala 109:76]
        writeStack_8_waitWFifoId <= _writeStack_8_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_33) begin // @[WriteStack.scala 115:15]
        writeStack_8_waitWFifoId <= _writeStack_8_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_8_waitWFifoId <= _GEN_680;
      end
    end else begin
      writeStack_8_waitWFifoId <= _GEN_680;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_35) begin // @[WriteStack.scala 109:76]
        writeStack_8_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_35) begin // @[WriteStack.scala 109:76]
        writeStack_8_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_8_validStatus <= _GEN_2449[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h8 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_8_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_8_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h8 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_8_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_59) begin // @[WriteStack.scala 233:15]
        writeStack_9_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_9_wvalid <= _GEN_297;
      end
    end else begin
      writeStack_9_wvalid <= _GEN_297;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h9 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_9_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_9_wstatus <= _GEN_2450[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h9 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_9_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_9_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h9 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_9_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_59) begin // @[WriteStack.scala 233:15]
        writeStack_9_entryFifoid <= _writeStack_9_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_681) begin // @[WriteStack.scala 240:15]
        writeStack_9_entryFifoid <= _writeStack_9_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_9_entryFifoid <= _GEN_1449;
      end
    end else begin
      writeStack_9_entryFifoid <= _GEN_1449;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_19 & _hasValid_T_28) begin // @[WriteStack.scala 151:84]
        writeStack_9_validFifoId <= _writeStack_9_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_19) begin // @[WriteStack.scala 154:65]
        writeStack_9_validFifoId <= _writeStack_9_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_9_validFifoId <= _GEN_1097;
      end
    end else begin
      writeStack_9_validFifoId <= _GEN_1097;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_39) begin // @[WriteStack.scala 109:76]
        writeStack_9_waitWFifoId <= _writeStack_9_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_37) begin // @[WriteStack.scala 115:15]
        writeStack_9_waitWFifoId <= _writeStack_9_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_9_waitWFifoId <= _GEN_681;
      end
    end else begin
      writeStack_9_waitWFifoId <= _GEN_681;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_39) begin // @[WriteStack.scala 109:76]
        writeStack_9_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_39) begin // @[WriteStack.scala 109:76]
        writeStack_9_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_9_validStatus <= _GEN_2451[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h9 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_9_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_9_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h9 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_9_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_65) begin // @[WriteStack.scala 233:15]
        writeStack_10_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_10_wvalid <= _GEN_298;
      end
    end else begin
      writeStack_10_wvalid <= _GEN_298;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'ha == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_10_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_10_wstatus <= _GEN_2452[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'ha == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_10_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_10_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'ha == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_10_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_65) begin // @[WriteStack.scala 233:15]
        writeStack_10_entryFifoid <= _writeStack_10_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_689) begin // @[WriteStack.scala 240:15]
        writeStack_10_entryFifoid <= _writeStack_10_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_10_entryFifoid <= _GEN_1450;
      end
    end else begin
      writeStack_10_entryFifoid <= _GEN_1450;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_21 & _hasValid_T_31) begin // @[WriteStack.scala 151:84]
        writeStack_10_validFifoId <= _writeStack_10_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_21) begin // @[WriteStack.scala 154:65]
        writeStack_10_validFifoId <= _writeStack_10_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_10_validFifoId <= _GEN_1098;
      end
    end else begin
      writeStack_10_validFifoId <= _GEN_1098;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_43) begin // @[WriteStack.scala 109:76]
        writeStack_10_waitWFifoId <= _writeStack_10_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_41) begin // @[WriteStack.scala 115:15]
        writeStack_10_waitWFifoId <= _writeStack_10_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_10_waitWFifoId <= _GEN_682;
      end
    end else begin
      writeStack_10_waitWFifoId <= _GEN_682;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_43) begin // @[WriteStack.scala 109:76]
        writeStack_10_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_43) begin // @[WriteStack.scala 109:76]
        writeStack_10_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_10_validStatus <= _GEN_2453[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'ha == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_10_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_10_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'ha == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_10_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_71) begin // @[WriteStack.scala 233:15]
        writeStack_11_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_11_wvalid <= _GEN_299;
      end
    end else begin
      writeStack_11_wvalid <= _GEN_299;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hb == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_11_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_11_wstatus <= _GEN_2454[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hb == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_11_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_11_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hb == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_11_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_71) begin // @[WriteStack.scala 233:15]
        writeStack_11_entryFifoid <= _writeStack_11_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_697) begin // @[WriteStack.scala 240:15]
        writeStack_11_entryFifoid <= _writeStack_11_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_11_entryFifoid <= _GEN_1451;
      end
    end else begin
      writeStack_11_entryFifoid <= _GEN_1451;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_23 & _hasValid_T_34) begin // @[WriteStack.scala 151:84]
        writeStack_11_validFifoId <= _writeStack_11_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_23) begin // @[WriteStack.scala 154:65]
        writeStack_11_validFifoId <= _writeStack_11_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_11_validFifoId <= _GEN_1099;
      end
    end else begin
      writeStack_11_validFifoId <= _GEN_1099;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_47) begin // @[WriteStack.scala 109:76]
        writeStack_11_waitWFifoId <= _writeStack_11_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_45) begin // @[WriteStack.scala 115:15]
        writeStack_11_waitWFifoId <= _writeStack_11_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_11_waitWFifoId <= _GEN_683;
      end
    end else begin
      writeStack_11_waitWFifoId <= _GEN_683;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_47) begin // @[WriteStack.scala 109:76]
        writeStack_11_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_47) begin // @[WriteStack.scala 109:76]
        writeStack_11_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_11_validStatus <= _GEN_2455[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hb == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_11_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_11_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hb == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_11_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_77) begin // @[WriteStack.scala 233:15]
        writeStack_12_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_12_wvalid <= _GEN_300;
      end
    end else begin
      writeStack_12_wvalid <= _GEN_300;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hc == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_12_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_12_wstatus <= _GEN_2456[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hc == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_12_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_12_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hc == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_12_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_77) begin // @[WriteStack.scala 233:15]
        writeStack_12_entryFifoid <= _writeStack_12_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_705) begin // @[WriteStack.scala 240:15]
        writeStack_12_entryFifoid <= _writeStack_12_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_12_entryFifoid <= _GEN_1452;
      end
    end else begin
      writeStack_12_entryFifoid <= _GEN_1452;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_25 & _hasValid_T_37) begin // @[WriteStack.scala 151:84]
        writeStack_12_validFifoId <= _writeStack_12_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_25) begin // @[WriteStack.scala 154:65]
        writeStack_12_validFifoId <= _writeStack_12_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_12_validFifoId <= _GEN_1100;
      end
    end else begin
      writeStack_12_validFifoId <= _GEN_1100;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_51) begin // @[WriteStack.scala 109:76]
        writeStack_12_waitWFifoId <= _writeStack_12_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_49) begin // @[WriteStack.scala 115:15]
        writeStack_12_waitWFifoId <= _writeStack_12_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_12_waitWFifoId <= _GEN_684;
      end
    end else begin
      writeStack_12_waitWFifoId <= _GEN_684;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_51) begin // @[WriteStack.scala 109:76]
        writeStack_12_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_51) begin // @[WriteStack.scala 109:76]
        writeStack_12_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_12_validStatus <= _GEN_2457[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hc == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_12_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_12_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hc == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_12_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_83) begin // @[WriteStack.scala 233:15]
        writeStack_13_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_13_wvalid <= _GEN_301;
      end
    end else begin
      writeStack_13_wvalid <= _GEN_301;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hd == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_13_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_13_wstatus <= _GEN_2458[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hd == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_13_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_13_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hd == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_13_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_83) begin // @[WriteStack.scala 233:15]
        writeStack_13_entryFifoid <= _writeStack_13_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_713) begin // @[WriteStack.scala 240:15]
        writeStack_13_entryFifoid <= _writeStack_13_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_13_entryFifoid <= _GEN_1453;
      end
    end else begin
      writeStack_13_entryFifoid <= _GEN_1453;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_27 & _hasValid_T_40) begin // @[WriteStack.scala 151:84]
        writeStack_13_validFifoId <= _writeStack_13_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_27) begin // @[WriteStack.scala 154:65]
        writeStack_13_validFifoId <= _writeStack_13_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_13_validFifoId <= _GEN_1101;
      end
    end else begin
      writeStack_13_validFifoId <= _GEN_1101;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_55) begin // @[WriteStack.scala 109:76]
        writeStack_13_waitWFifoId <= _writeStack_13_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_53) begin // @[WriteStack.scala 115:15]
        writeStack_13_waitWFifoId <= _writeStack_13_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_13_waitWFifoId <= _GEN_685;
      end
    end else begin
      writeStack_13_waitWFifoId <= _GEN_685;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_55) begin // @[WriteStack.scala 109:76]
        writeStack_13_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_55) begin // @[WriteStack.scala 109:76]
        writeStack_13_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_13_validStatus <= _GEN_2459[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hd == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_13_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_13_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hd == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_13_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_89) begin // @[WriteStack.scala 233:15]
        writeStack_14_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_14_wvalid <= _GEN_302;
      end
    end else begin
      writeStack_14_wvalid <= _GEN_302;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'he == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_14_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_14_wstatus <= _GEN_2460[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'he == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_14_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_14_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'he == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_14_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_89) begin // @[WriteStack.scala 233:15]
        writeStack_14_entryFifoid <= _writeStack_14_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_721) begin // @[WriteStack.scala 240:15]
        writeStack_14_entryFifoid <= _writeStack_14_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_14_entryFifoid <= _GEN_1454;
      end
    end else begin
      writeStack_14_entryFifoid <= _GEN_1454;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_29 & _hasValid_T_43) begin // @[WriteStack.scala 151:84]
        writeStack_14_validFifoId <= _writeStack_14_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_29) begin // @[WriteStack.scala 154:65]
        writeStack_14_validFifoId <= _writeStack_14_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_14_validFifoId <= _GEN_1102;
      end
    end else begin
      writeStack_14_validFifoId <= _GEN_1102;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_59) begin // @[WriteStack.scala 109:76]
        writeStack_14_waitWFifoId <= _writeStack_14_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_57) begin // @[WriteStack.scala 115:15]
        writeStack_14_waitWFifoId <= _writeStack_14_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_14_waitWFifoId <= _GEN_686;
      end
    end else begin
      writeStack_14_waitWFifoId <= _GEN_686;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_59) begin // @[WriteStack.scala 109:76]
        writeStack_14_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_59) begin // @[WriteStack.scala 109:76]
        writeStack_14_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_14_validStatus <= _GEN_2461[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'he == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_14_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_14_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'he == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_14_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_95) begin // @[WriteStack.scala 233:15]
        writeStack_15_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_15_wvalid <= _GEN_303;
      end
    end else begin
      writeStack_15_wvalid <= _GEN_303;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hf == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_15_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_15_wstatus <= _GEN_2462[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hf == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_15_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_15_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hf == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_15_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_95) begin // @[WriteStack.scala 233:15]
        writeStack_15_entryFifoid <= _writeStack_15_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_729) begin // @[WriteStack.scala 240:15]
        writeStack_15_entryFifoid <= _writeStack_15_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_15_entryFifoid <= _GEN_1455;
      end
    end else begin
      writeStack_15_entryFifoid <= _GEN_1455;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_31 & _hasValid_T_46) begin // @[WriteStack.scala 151:84]
        writeStack_15_validFifoId <= _writeStack_15_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_31) begin // @[WriteStack.scala 154:65]
        writeStack_15_validFifoId <= _writeStack_15_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_15_validFifoId <= _GEN_1103;
      end
    end else begin
      writeStack_15_validFifoId <= _GEN_1103;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_63) begin // @[WriteStack.scala 109:76]
        writeStack_15_waitWFifoId <= _writeStack_15_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_61) begin // @[WriteStack.scala 115:15]
        writeStack_15_waitWFifoId <= _writeStack_15_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_15_waitWFifoId <= _GEN_687;
      end
    end else begin
      writeStack_15_waitWFifoId <= _GEN_687;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_63) begin // @[WriteStack.scala 109:76]
        writeStack_15_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_63) begin // @[WriteStack.scala 109:76]
        writeStack_15_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_15_validStatus <= _GEN_2463[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hf == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_15_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_15_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'hf == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_15_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_101) begin // @[WriteStack.scala 233:15]
        writeStack_16_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_16_wvalid <= _GEN_304;
      end
    end else begin
      writeStack_16_wvalid <= _GEN_304;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h10 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_16_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_16_wstatus <= _GEN_2464[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h10 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_16_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_16_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h10 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_16_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_101) begin // @[WriteStack.scala 233:15]
        writeStack_16_entryFifoid <= _writeStack_16_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_737) begin // @[WriteStack.scala 240:15]
        writeStack_16_entryFifoid <= _writeStack_16_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_16_entryFifoid <= _GEN_1456;
      end
    end else begin
      writeStack_16_entryFifoid <= _GEN_1456;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_33 & _hasValid_T_49) begin // @[WriteStack.scala 151:84]
        writeStack_16_validFifoId <= _writeStack_16_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_33) begin // @[WriteStack.scala 154:65]
        writeStack_16_validFifoId <= _writeStack_16_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_16_validFifoId <= _GEN_1104;
      end
    end else begin
      writeStack_16_validFifoId <= _GEN_1104;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_67) begin // @[WriteStack.scala 109:76]
        writeStack_16_waitWFifoId <= _writeStack_16_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_65) begin // @[WriteStack.scala 115:15]
        writeStack_16_waitWFifoId <= _writeStack_16_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_16_waitWFifoId <= _GEN_688;
      end
    end else begin
      writeStack_16_waitWFifoId <= _GEN_688;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_67) begin // @[WriteStack.scala 109:76]
        writeStack_16_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_67) begin // @[WriteStack.scala 109:76]
        writeStack_16_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_16_validStatus <= _GEN_2465[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h10 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_16_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_16_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h10 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_16_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_107) begin // @[WriteStack.scala 233:15]
        writeStack_17_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_17_wvalid <= _GEN_305;
      end
    end else begin
      writeStack_17_wvalid <= _GEN_305;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h11 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_17_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_17_wstatus <= _GEN_2466[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h11 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_17_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_17_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h11 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_17_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_107) begin // @[WriteStack.scala 233:15]
        writeStack_17_entryFifoid <= _writeStack_17_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_745) begin // @[WriteStack.scala 240:15]
        writeStack_17_entryFifoid <= _writeStack_17_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_17_entryFifoid <= _GEN_1457;
      end
    end else begin
      writeStack_17_entryFifoid <= _GEN_1457;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_35 & _hasValid_T_52) begin // @[WriteStack.scala 151:84]
        writeStack_17_validFifoId <= _writeStack_17_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_35) begin // @[WriteStack.scala 154:65]
        writeStack_17_validFifoId <= _writeStack_17_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_17_validFifoId <= _GEN_1105;
      end
    end else begin
      writeStack_17_validFifoId <= _GEN_1105;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_71) begin // @[WriteStack.scala 109:76]
        writeStack_17_waitWFifoId <= _writeStack_17_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_69) begin // @[WriteStack.scala 115:15]
        writeStack_17_waitWFifoId <= _writeStack_17_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_17_waitWFifoId <= _GEN_689;
      end
    end else begin
      writeStack_17_waitWFifoId <= _GEN_689;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_71) begin // @[WriteStack.scala 109:76]
        writeStack_17_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_71) begin // @[WriteStack.scala 109:76]
        writeStack_17_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_17_validStatus <= _GEN_2467[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h11 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_17_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_17_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h11 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_17_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_113) begin // @[WriteStack.scala 233:15]
        writeStack_18_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_18_wvalid <= _GEN_306;
      end
    end else begin
      writeStack_18_wvalid <= _GEN_306;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h12 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_18_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_18_wstatus <= _GEN_2468[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h12 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_18_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_18_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h12 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_18_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_113) begin // @[WriteStack.scala 233:15]
        writeStack_18_entryFifoid <= _writeStack_18_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_753) begin // @[WriteStack.scala 240:15]
        writeStack_18_entryFifoid <= _writeStack_18_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_18_entryFifoid <= _GEN_1458;
      end
    end else begin
      writeStack_18_entryFifoid <= _GEN_1458;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_37 & _hasValid_T_55) begin // @[WriteStack.scala 151:84]
        writeStack_18_validFifoId <= _writeStack_18_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_37) begin // @[WriteStack.scala 154:65]
        writeStack_18_validFifoId <= _writeStack_18_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_18_validFifoId <= _GEN_1106;
      end
    end else begin
      writeStack_18_validFifoId <= _GEN_1106;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_75) begin // @[WriteStack.scala 109:76]
        writeStack_18_waitWFifoId <= _writeStack_18_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_73) begin // @[WriteStack.scala 115:15]
        writeStack_18_waitWFifoId <= _writeStack_18_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_18_waitWFifoId <= _GEN_690;
      end
    end else begin
      writeStack_18_waitWFifoId <= _GEN_690;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_75) begin // @[WriteStack.scala 109:76]
        writeStack_18_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_75) begin // @[WriteStack.scala 109:76]
        writeStack_18_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_18_validStatus <= _GEN_2469[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h12 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_18_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_18_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h12 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_18_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_119) begin // @[WriteStack.scala 233:15]
        writeStack_19_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_19_wvalid <= _GEN_307;
      end
    end else begin
      writeStack_19_wvalid <= _GEN_307;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h13 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_19_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_19_wstatus <= _GEN_2470[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h13 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_19_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_19_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h13 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_19_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_119) begin // @[WriteStack.scala 233:15]
        writeStack_19_entryFifoid <= _writeStack_19_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_761) begin // @[WriteStack.scala 240:15]
        writeStack_19_entryFifoid <= _writeStack_19_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_19_entryFifoid <= _GEN_1459;
      end
    end else begin
      writeStack_19_entryFifoid <= _GEN_1459;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_39 & _hasValid_T_58) begin // @[WriteStack.scala 151:84]
        writeStack_19_validFifoId <= _writeStack_19_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_39) begin // @[WriteStack.scala 154:65]
        writeStack_19_validFifoId <= _writeStack_19_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_19_validFifoId <= _GEN_1107;
      end
    end else begin
      writeStack_19_validFifoId <= _GEN_1107;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_79) begin // @[WriteStack.scala 109:76]
        writeStack_19_waitWFifoId <= _writeStack_19_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_77) begin // @[WriteStack.scala 115:15]
        writeStack_19_waitWFifoId <= _writeStack_19_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_19_waitWFifoId <= _GEN_691;
      end
    end else begin
      writeStack_19_waitWFifoId <= _GEN_691;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_79) begin // @[WriteStack.scala 109:76]
        writeStack_19_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_79) begin // @[WriteStack.scala 109:76]
        writeStack_19_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_19_validStatus <= _GEN_2471[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h13 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_19_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_19_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h13 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_19_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_125) begin // @[WriteStack.scala 233:15]
        writeStack_20_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_20_wvalid <= _GEN_308;
      end
    end else begin
      writeStack_20_wvalid <= _GEN_308;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h14 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_20_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_20_wstatus <= _GEN_2472[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h14 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_20_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_20_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h14 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_20_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_125) begin // @[WriteStack.scala 233:15]
        writeStack_20_entryFifoid <= _writeStack_20_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_769) begin // @[WriteStack.scala 240:15]
        writeStack_20_entryFifoid <= _writeStack_20_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_20_entryFifoid <= _GEN_1460;
      end
    end else begin
      writeStack_20_entryFifoid <= _GEN_1460;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_41 & _hasValid_T_61) begin // @[WriteStack.scala 151:84]
        writeStack_20_validFifoId <= _writeStack_20_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_41) begin // @[WriteStack.scala 154:65]
        writeStack_20_validFifoId <= _writeStack_20_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_20_validFifoId <= _GEN_1108;
      end
    end else begin
      writeStack_20_validFifoId <= _GEN_1108;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_83) begin // @[WriteStack.scala 109:76]
        writeStack_20_waitWFifoId <= _writeStack_20_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_81) begin // @[WriteStack.scala 115:15]
        writeStack_20_waitWFifoId <= _writeStack_20_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_20_waitWFifoId <= _GEN_692;
      end
    end else begin
      writeStack_20_waitWFifoId <= _GEN_692;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_83) begin // @[WriteStack.scala 109:76]
        writeStack_20_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_83) begin // @[WriteStack.scala 109:76]
        writeStack_20_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_20_validStatus <= _GEN_2473[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h14 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_20_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_20_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h14 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_20_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_131) begin // @[WriteStack.scala 233:15]
        writeStack_21_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_21_wvalid <= _GEN_309;
      end
    end else begin
      writeStack_21_wvalid <= _GEN_309;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h15 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_21_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_21_wstatus <= _GEN_2474[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h15 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_21_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_21_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h15 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_21_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_131) begin // @[WriteStack.scala 233:15]
        writeStack_21_entryFifoid <= _writeStack_21_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_777) begin // @[WriteStack.scala 240:15]
        writeStack_21_entryFifoid <= _writeStack_21_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_21_entryFifoid <= _GEN_1461;
      end
    end else begin
      writeStack_21_entryFifoid <= _GEN_1461;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_43 & _hasValid_T_64) begin // @[WriteStack.scala 151:84]
        writeStack_21_validFifoId <= _writeStack_21_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_43) begin // @[WriteStack.scala 154:65]
        writeStack_21_validFifoId <= _writeStack_21_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_21_validFifoId <= _GEN_1109;
      end
    end else begin
      writeStack_21_validFifoId <= _GEN_1109;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_87) begin // @[WriteStack.scala 109:76]
        writeStack_21_waitWFifoId <= _writeStack_21_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_85) begin // @[WriteStack.scala 115:15]
        writeStack_21_waitWFifoId <= _writeStack_21_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_21_waitWFifoId <= _GEN_693;
      end
    end else begin
      writeStack_21_waitWFifoId <= _GEN_693;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_87) begin // @[WriteStack.scala 109:76]
        writeStack_21_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_87) begin // @[WriteStack.scala 109:76]
        writeStack_21_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_21_validStatus <= _GEN_2475[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h15 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_21_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_21_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h15 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_21_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_137) begin // @[WriteStack.scala 233:15]
        writeStack_22_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_22_wvalid <= _GEN_310;
      end
    end else begin
      writeStack_22_wvalid <= _GEN_310;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h16 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_22_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_22_wstatus <= _GEN_2476[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h16 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_22_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_22_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h16 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_22_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_137) begin // @[WriteStack.scala 233:15]
        writeStack_22_entryFifoid <= _writeStack_22_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_785) begin // @[WriteStack.scala 240:15]
        writeStack_22_entryFifoid <= _writeStack_22_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_22_entryFifoid <= _GEN_1462;
      end
    end else begin
      writeStack_22_entryFifoid <= _GEN_1462;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_45 & _hasValid_T_67) begin // @[WriteStack.scala 151:84]
        writeStack_22_validFifoId <= _writeStack_22_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_45) begin // @[WriteStack.scala 154:65]
        writeStack_22_validFifoId <= _writeStack_22_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_22_validFifoId <= _GEN_1110;
      end
    end else begin
      writeStack_22_validFifoId <= _GEN_1110;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_91) begin // @[WriteStack.scala 109:76]
        writeStack_22_waitWFifoId <= _writeStack_22_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_89) begin // @[WriteStack.scala 115:15]
        writeStack_22_waitWFifoId <= _writeStack_22_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_22_waitWFifoId <= _GEN_694;
      end
    end else begin
      writeStack_22_waitWFifoId <= _GEN_694;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_91) begin // @[WriteStack.scala 109:76]
        writeStack_22_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_91) begin // @[WriteStack.scala 109:76]
        writeStack_22_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_22_validStatus <= _GEN_2477[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h16 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_22_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_22_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h16 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_22_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_143) begin // @[WriteStack.scala 233:15]
        writeStack_23_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_23_wvalid <= _GEN_311;
      end
    end else begin
      writeStack_23_wvalid <= _GEN_311;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h17 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_23_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_23_wstatus <= _GEN_2478[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h17 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_23_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_23_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h17 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_23_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_143) begin // @[WriteStack.scala 233:15]
        writeStack_23_entryFifoid <= _writeStack_23_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_793) begin // @[WriteStack.scala 240:15]
        writeStack_23_entryFifoid <= _writeStack_23_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_23_entryFifoid <= _GEN_1463;
      end
    end else begin
      writeStack_23_entryFifoid <= _GEN_1463;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_47 & _hasValid_T_70) begin // @[WriteStack.scala 151:84]
        writeStack_23_validFifoId <= _writeStack_23_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_47) begin // @[WriteStack.scala 154:65]
        writeStack_23_validFifoId <= _writeStack_23_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_23_validFifoId <= _GEN_1111;
      end
    end else begin
      writeStack_23_validFifoId <= _GEN_1111;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_95) begin // @[WriteStack.scala 109:76]
        writeStack_23_waitWFifoId <= _writeStack_23_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_93) begin // @[WriteStack.scala 115:15]
        writeStack_23_waitWFifoId <= _writeStack_23_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_23_waitWFifoId <= _GEN_695;
      end
    end else begin
      writeStack_23_waitWFifoId <= _GEN_695;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_95) begin // @[WriteStack.scala 109:76]
        writeStack_23_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_95) begin // @[WriteStack.scala 109:76]
        writeStack_23_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_23_validStatus <= _GEN_2479[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h17 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_23_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_23_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h17 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_23_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_149) begin // @[WriteStack.scala 233:15]
        writeStack_24_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_24_wvalid <= _GEN_312;
      end
    end else begin
      writeStack_24_wvalid <= _GEN_312;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h18 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_24_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_24_wstatus <= _GEN_2480[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h18 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_24_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_24_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h18 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_24_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_149) begin // @[WriteStack.scala 233:15]
        writeStack_24_entryFifoid <= _writeStack_24_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_801) begin // @[WriteStack.scala 240:15]
        writeStack_24_entryFifoid <= _writeStack_24_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_24_entryFifoid <= _GEN_1464;
      end
    end else begin
      writeStack_24_entryFifoid <= _GEN_1464;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_49 & _hasValid_T_73) begin // @[WriteStack.scala 151:84]
        writeStack_24_validFifoId <= _writeStack_24_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_49) begin // @[WriteStack.scala 154:65]
        writeStack_24_validFifoId <= _writeStack_24_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_24_validFifoId <= _GEN_1112;
      end
    end else begin
      writeStack_24_validFifoId <= _GEN_1112;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_99) begin // @[WriteStack.scala 109:76]
        writeStack_24_waitWFifoId <= _writeStack_24_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_97) begin // @[WriteStack.scala 115:15]
        writeStack_24_waitWFifoId <= _writeStack_24_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_24_waitWFifoId <= _GEN_696;
      end
    end else begin
      writeStack_24_waitWFifoId <= _GEN_696;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_99) begin // @[WriteStack.scala 109:76]
        writeStack_24_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_99) begin // @[WriteStack.scala 109:76]
        writeStack_24_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_24_validStatus <= _GEN_2481[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h18 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_24_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_24_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h18 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_24_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_155) begin // @[WriteStack.scala 233:15]
        writeStack_25_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_25_wvalid <= _GEN_313;
      end
    end else begin
      writeStack_25_wvalid <= _GEN_313;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h19 == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_25_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_25_wstatus <= _GEN_2482[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h19 == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_25_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_25_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h19 == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_25_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_155) begin // @[WriteStack.scala 233:15]
        writeStack_25_entryFifoid <= _writeStack_25_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_809) begin // @[WriteStack.scala 240:15]
        writeStack_25_entryFifoid <= _writeStack_25_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_25_entryFifoid <= _GEN_1465;
      end
    end else begin
      writeStack_25_entryFifoid <= _GEN_1465;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_51 & _hasValid_T_76) begin // @[WriteStack.scala 151:84]
        writeStack_25_validFifoId <= _writeStack_25_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_51) begin // @[WriteStack.scala 154:65]
        writeStack_25_validFifoId <= _writeStack_25_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_25_validFifoId <= _GEN_1113;
      end
    end else begin
      writeStack_25_validFifoId <= _GEN_1113;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_103) begin // @[WriteStack.scala 109:76]
        writeStack_25_waitWFifoId <= _writeStack_25_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_101) begin // @[WriteStack.scala 115:15]
        writeStack_25_waitWFifoId <= _writeStack_25_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_25_waitWFifoId <= _GEN_697;
      end
    end else begin
      writeStack_25_waitWFifoId <= _GEN_697;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_103) begin // @[WriteStack.scala 109:76]
        writeStack_25_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_103) begin // @[WriteStack.scala 109:76]
        writeStack_25_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_25_validStatus <= _GEN_2483[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h19 == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_25_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_25_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h19 == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_25_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_161) begin // @[WriteStack.scala 233:15]
        writeStack_26_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_26_wvalid <= _GEN_314;
      end
    end else begin
      writeStack_26_wvalid <= _GEN_314;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1a == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_26_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_26_wstatus <= _GEN_2484[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1a == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_26_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_26_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1a == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_26_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_161) begin // @[WriteStack.scala 233:15]
        writeStack_26_entryFifoid <= _writeStack_26_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_817) begin // @[WriteStack.scala 240:15]
        writeStack_26_entryFifoid <= _writeStack_26_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_26_entryFifoid <= _GEN_1466;
      end
    end else begin
      writeStack_26_entryFifoid <= _GEN_1466;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_53 & _hasValid_T_79) begin // @[WriteStack.scala 151:84]
        writeStack_26_validFifoId <= _writeStack_26_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_53) begin // @[WriteStack.scala 154:65]
        writeStack_26_validFifoId <= _writeStack_26_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_26_validFifoId <= _GEN_1114;
      end
    end else begin
      writeStack_26_validFifoId <= _GEN_1114;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_107) begin // @[WriteStack.scala 109:76]
        writeStack_26_waitWFifoId <= _writeStack_26_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_105) begin // @[WriteStack.scala 115:15]
        writeStack_26_waitWFifoId <= _writeStack_26_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_26_waitWFifoId <= _GEN_698;
      end
    end else begin
      writeStack_26_waitWFifoId <= _GEN_698;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_107) begin // @[WriteStack.scala 109:76]
        writeStack_26_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_107) begin // @[WriteStack.scala 109:76]
        writeStack_26_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_26_validStatus <= _GEN_2485[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1a == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_26_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_26_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1a == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_26_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_167) begin // @[WriteStack.scala 233:15]
        writeStack_27_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_27_wvalid <= _GEN_315;
      end
    end else begin
      writeStack_27_wvalid <= _GEN_315;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1b == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_27_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_27_wstatus <= _GEN_2486[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1b == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_27_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_27_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1b == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_27_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_167) begin // @[WriteStack.scala 233:15]
        writeStack_27_entryFifoid <= _writeStack_27_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_825) begin // @[WriteStack.scala 240:15]
        writeStack_27_entryFifoid <= _writeStack_27_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_27_entryFifoid <= _GEN_1467;
      end
    end else begin
      writeStack_27_entryFifoid <= _GEN_1467;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_55 & _hasValid_T_82) begin // @[WriteStack.scala 151:84]
        writeStack_27_validFifoId <= _writeStack_27_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_55) begin // @[WriteStack.scala 154:65]
        writeStack_27_validFifoId <= _writeStack_27_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_27_validFifoId <= _GEN_1115;
      end
    end else begin
      writeStack_27_validFifoId <= _GEN_1115;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_111) begin // @[WriteStack.scala 109:76]
        writeStack_27_waitWFifoId <= _writeStack_27_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_109) begin // @[WriteStack.scala 115:15]
        writeStack_27_waitWFifoId <= _writeStack_27_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_27_waitWFifoId <= _GEN_699;
      end
    end else begin
      writeStack_27_waitWFifoId <= _GEN_699;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_111) begin // @[WriteStack.scala 109:76]
        writeStack_27_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_111) begin // @[WriteStack.scala 109:76]
        writeStack_27_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_27_validStatus <= _GEN_2487[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1b == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_27_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_27_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1b == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_27_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_173) begin // @[WriteStack.scala 233:15]
        writeStack_28_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_28_wvalid <= _GEN_316;
      end
    end else begin
      writeStack_28_wvalid <= _GEN_316;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1c == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_28_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_28_wstatus <= _GEN_2488[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1c == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_28_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_28_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1c == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_28_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_173) begin // @[WriteStack.scala 233:15]
        writeStack_28_entryFifoid <= _writeStack_28_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_833) begin // @[WriteStack.scala 240:15]
        writeStack_28_entryFifoid <= _writeStack_28_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_28_entryFifoid <= _GEN_1468;
      end
    end else begin
      writeStack_28_entryFifoid <= _GEN_1468;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_57 & _hasValid_T_85) begin // @[WriteStack.scala 151:84]
        writeStack_28_validFifoId <= _writeStack_28_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_57) begin // @[WriteStack.scala 154:65]
        writeStack_28_validFifoId <= _writeStack_28_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_28_validFifoId <= _GEN_1116;
      end
    end else begin
      writeStack_28_validFifoId <= _GEN_1116;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_115) begin // @[WriteStack.scala 109:76]
        writeStack_28_waitWFifoId <= _writeStack_28_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_113) begin // @[WriteStack.scala 115:15]
        writeStack_28_waitWFifoId <= _writeStack_28_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_28_waitWFifoId <= _GEN_700;
      end
    end else begin
      writeStack_28_waitWFifoId <= _GEN_700;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_115) begin // @[WriteStack.scala 109:76]
        writeStack_28_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_115) begin // @[WriteStack.scala 109:76]
        writeStack_28_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_28_validStatus <= _GEN_2489[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1c == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_28_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_28_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1c == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_28_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_179) begin // @[WriteStack.scala 233:15]
        writeStack_29_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_29_wvalid <= _GEN_317;
      end
    end else begin
      writeStack_29_wvalid <= _GEN_317;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1d == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_29_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_29_wstatus <= _GEN_2490[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1d == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_29_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_29_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1d == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_29_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_179) begin // @[WriteStack.scala 233:15]
        writeStack_29_entryFifoid <= _writeStack_29_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_841) begin // @[WriteStack.scala 240:15]
        writeStack_29_entryFifoid <= _writeStack_29_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_29_entryFifoid <= _GEN_1469;
      end
    end else begin
      writeStack_29_entryFifoid <= _GEN_1469;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_59 & _hasValid_T_88) begin // @[WriteStack.scala 151:84]
        writeStack_29_validFifoId <= _writeStack_29_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_59) begin // @[WriteStack.scala 154:65]
        writeStack_29_validFifoId <= _writeStack_29_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_29_validFifoId <= _GEN_1117;
      end
    end else begin
      writeStack_29_validFifoId <= _GEN_1117;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_119) begin // @[WriteStack.scala 109:76]
        writeStack_29_waitWFifoId <= _writeStack_29_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_117) begin // @[WriteStack.scala 115:15]
        writeStack_29_waitWFifoId <= _writeStack_29_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_29_waitWFifoId <= _GEN_701;
      end
    end else begin
      writeStack_29_waitWFifoId <= _GEN_701;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_119) begin // @[WriteStack.scala 109:76]
        writeStack_29_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_119) begin // @[WriteStack.scala 109:76]
        writeStack_29_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_29_validStatus <= _GEN_2491[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1d == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_29_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_29_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1d == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_29_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_185) begin // @[WriteStack.scala 233:15]
        writeStack_30_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_30_wvalid <= _GEN_318;
      end
    end else begin
      writeStack_30_wvalid <= _GEN_318;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1e == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_30_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_30_wstatus <= _GEN_2492[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1e == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_30_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_30_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1e == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_30_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_185) begin // @[WriteStack.scala 233:15]
        writeStack_30_entryFifoid <= _writeStack_30_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_849) begin // @[WriteStack.scala 240:15]
        writeStack_30_entryFifoid <= _writeStack_30_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_30_entryFifoid <= _GEN_1470;
      end
    end else begin
      writeStack_30_entryFifoid <= _GEN_1470;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_61 & _hasValid_T_91) begin // @[WriteStack.scala 151:84]
        writeStack_30_validFifoId <= _writeStack_30_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_61) begin // @[WriteStack.scala 154:65]
        writeStack_30_validFifoId <= _writeStack_30_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_30_validFifoId <= _GEN_1118;
      end
    end else begin
      writeStack_30_validFifoId <= _GEN_1118;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_123) begin // @[WriteStack.scala 109:76]
        writeStack_30_waitWFifoId <= _writeStack_30_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_121) begin // @[WriteStack.scala 115:15]
        writeStack_30_waitWFifoId <= _writeStack_30_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_30_waitWFifoId <= _GEN_702;
      end
    end else begin
      writeStack_30_waitWFifoId <= _GEN_702;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_123) begin // @[WriteStack.scala 109:76]
        writeStack_30_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_123) begin // @[WriteStack.scala 109:76]
        writeStack_30_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_30_validStatus <= _GEN_2493[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1e == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_30_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_30_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1e == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_30_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_wvalid <= 1'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_191) begin // @[WriteStack.scala 233:15]
        writeStack_31_wvalid <= 1'h0; // @[WriteStack.scala 236:28]
      end else begin
        writeStack_31_wvalid <= _GEN_319;
      end
    end else begin
      writeStack_31_wvalid <= _GEN_319;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_waddr <= 35'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1f == idxInsert) begin // @[WriteStack.scala 74:17]
        writeStack_31_waddr <= io_axiWriteReq_in_aw_bits_addr; // @[WriteStack.scala 74:17]
      end
    end
    writeStack_31_wstatus <= _GEN_2494[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_entryid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1f == idxInsert) begin // @[WriteStack.scala 81:19]
        if (alloc) begin // @[WriteStack.scala 68:22]
          writeStack_31_entryid <= _idxInsert_T_62;
        end else begin
          writeStack_31_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_awid <= 14'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1f == idxInsert) begin // @[WriteStack.scala 80:16]
        writeStack_31_awid <= io_axiWriteReq_in_aw_bits_id; // @[WriteStack.scala 80:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_entryFifoid <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_402) begin // @[WriteStack.scala 229:3]
      if (_canMenW_T_191) begin // @[WriteStack.scala 233:15]
        writeStack_31_entryFifoid <= _writeStack_31_entryFifoid_T_1; // @[WriteStack.scala 238:33]
      end else if (_T_857) begin // @[WriteStack.scala 240:15]
        writeStack_31_entryFifoid <= _writeStack_31_entryFifoid_T_1; // @[WriteStack.scala 241:33]
      end else begin
        writeStack_31_entryFifoid <= _GEN_1471;
      end
    end else begin
      writeStack_31_entryFifoid <= _GEN_1471;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_validFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_201) begin // @[WriteStack.scala 148:5]
      if (_writeStack_validFifoId_T_63 & _hasValid_T_94) begin // @[WriteStack.scala 151:84]
        writeStack_31_validFifoId <= _writeStack_31_validFifoId_T_1; // @[WriteStack.scala 153:29]
      end else if (_writeStack_validFifoId_T_63) begin // @[WriteStack.scala 154:65]
        writeStack_31_validFifoId <= _writeStack_31_validFifoId_T_1; // @[WriteStack.scala 155:29]
      end else begin
        writeStack_31_validFifoId <= _GEN_1119;
      end
    end else begin
      writeStack_31_validFifoId <= _GEN_1119;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_waitWFifoId <= 5'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_127) begin // @[WriteStack.scala 109:76]
        writeStack_31_waitWFifoId <= _writeStack_31_waitWFifoId_T_1; // @[WriteStack.scala 113:31]
      end else if (_canW_T_125) begin // @[WriteStack.scala 115:15]
        writeStack_31_waitWFifoId <= _writeStack_31_waitWFifoId_T_1; // @[WriteStack.scala 116:31]
      end else begin
        writeStack_31_waitWFifoId <= _GEN_703;
      end
    end else begin
      writeStack_31_waitWFifoId <= _GEN_703;
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_data <= 256'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_127) begin // @[WriteStack.scala 109:76]
        writeStack_31_data <= io_axiWriteReq_in_w_bits_data; // @[WriteStack.scala 110:24]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_mask <= 32'h0; // @[WriteStack.scala 56:27]
    end else if (_T_1) begin // @[WriteStack.scala 106:5]
      if (_canW_T_127) begin // @[WriteStack.scala 109:76]
        writeStack_31_mask <= io_axiWriteReq_in_w_bits_strb; // @[WriteStack.scala 111:24]
      end
    end
    writeStack_31_validStatus <= _GEN_2495[1:0]; // @[WriteStack.scala 56:{27,27}]
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_size <= 3'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1f == idxInsert) begin // @[WriteStack.scala 78:16]
        writeStack_31_size <= io_axiWriteReq_in_aw_bits_size; // @[WriteStack.scala 78:16]
      end
    end
    if (reset) begin // @[WriteStack.scala 56:27]
      writeStack_31_len <= 8'h0; // @[WriteStack.scala 56:27]
    end else if (alloc) begin // @[WriteStack.scala 70:14]
      if (5'h1f == idxInsert) begin // @[WriteStack.scala 79:15]
        writeStack_31_len <= io_axiWriteReq_in_aw_bits_len; // @[WriteStack.scala 79:15]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  writeStack_0_wvalid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  writeStack_0_waddr = _RAND_1[34:0];
  _RAND_2 = {1{`RANDOM}};
  writeStack_0_wstatus = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  writeStack_0_entryid = _RAND_3[4:0];
  _RAND_4 = {1{`RANDOM}};
  writeStack_0_awid = _RAND_4[13:0];
  _RAND_5 = {1{`RANDOM}};
  writeStack_0_entryFifoid = _RAND_5[4:0];
  _RAND_6 = {1{`RANDOM}};
  writeStack_0_validFifoId = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  writeStack_0_waitWFifoId = _RAND_7[4:0];
  _RAND_8 = {8{`RANDOM}};
  writeStack_0_data = _RAND_8[255:0];
  _RAND_9 = {1{`RANDOM}};
  writeStack_0_mask = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  writeStack_0_validStatus = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  writeStack_0_size = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  writeStack_0_len = _RAND_12[7:0];
  _RAND_13 = {1{`RANDOM}};
  writeStack_1_wvalid = _RAND_13[0:0];
  _RAND_14 = {2{`RANDOM}};
  writeStack_1_waddr = _RAND_14[34:0];
  _RAND_15 = {1{`RANDOM}};
  writeStack_1_wstatus = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  writeStack_1_entryid = _RAND_16[4:0];
  _RAND_17 = {1{`RANDOM}};
  writeStack_1_awid = _RAND_17[13:0];
  _RAND_18 = {1{`RANDOM}};
  writeStack_1_entryFifoid = _RAND_18[4:0];
  _RAND_19 = {1{`RANDOM}};
  writeStack_1_validFifoId = _RAND_19[4:0];
  _RAND_20 = {1{`RANDOM}};
  writeStack_1_waitWFifoId = _RAND_20[4:0];
  _RAND_21 = {8{`RANDOM}};
  writeStack_1_data = _RAND_21[255:0];
  _RAND_22 = {1{`RANDOM}};
  writeStack_1_mask = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  writeStack_1_validStatus = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  writeStack_1_size = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  writeStack_1_len = _RAND_25[7:0];
  _RAND_26 = {1{`RANDOM}};
  writeStack_2_wvalid = _RAND_26[0:0];
  _RAND_27 = {2{`RANDOM}};
  writeStack_2_waddr = _RAND_27[34:0];
  _RAND_28 = {1{`RANDOM}};
  writeStack_2_wstatus = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  writeStack_2_entryid = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  writeStack_2_awid = _RAND_30[13:0];
  _RAND_31 = {1{`RANDOM}};
  writeStack_2_entryFifoid = _RAND_31[4:0];
  _RAND_32 = {1{`RANDOM}};
  writeStack_2_validFifoId = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  writeStack_2_waitWFifoId = _RAND_33[4:0];
  _RAND_34 = {8{`RANDOM}};
  writeStack_2_data = _RAND_34[255:0];
  _RAND_35 = {1{`RANDOM}};
  writeStack_2_mask = _RAND_35[31:0];
  _RAND_36 = {1{`RANDOM}};
  writeStack_2_validStatus = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  writeStack_2_size = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  writeStack_2_len = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  writeStack_3_wvalid = _RAND_39[0:0];
  _RAND_40 = {2{`RANDOM}};
  writeStack_3_waddr = _RAND_40[34:0];
  _RAND_41 = {1{`RANDOM}};
  writeStack_3_wstatus = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  writeStack_3_entryid = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  writeStack_3_awid = _RAND_43[13:0];
  _RAND_44 = {1{`RANDOM}};
  writeStack_3_entryFifoid = _RAND_44[4:0];
  _RAND_45 = {1{`RANDOM}};
  writeStack_3_validFifoId = _RAND_45[4:0];
  _RAND_46 = {1{`RANDOM}};
  writeStack_3_waitWFifoId = _RAND_46[4:0];
  _RAND_47 = {8{`RANDOM}};
  writeStack_3_data = _RAND_47[255:0];
  _RAND_48 = {1{`RANDOM}};
  writeStack_3_mask = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  writeStack_3_validStatus = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  writeStack_3_size = _RAND_50[2:0];
  _RAND_51 = {1{`RANDOM}};
  writeStack_3_len = _RAND_51[7:0];
  _RAND_52 = {1{`RANDOM}};
  writeStack_4_wvalid = _RAND_52[0:0];
  _RAND_53 = {2{`RANDOM}};
  writeStack_4_waddr = _RAND_53[34:0];
  _RAND_54 = {1{`RANDOM}};
  writeStack_4_wstatus = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  writeStack_4_entryid = _RAND_55[4:0];
  _RAND_56 = {1{`RANDOM}};
  writeStack_4_awid = _RAND_56[13:0];
  _RAND_57 = {1{`RANDOM}};
  writeStack_4_entryFifoid = _RAND_57[4:0];
  _RAND_58 = {1{`RANDOM}};
  writeStack_4_validFifoId = _RAND_58[4:0];
  _RAND_59 = {1{`RANDOM}};
  writeStack_4_waitWFifoId = _RAND_59[4:0];
  _RAND_60 = {8{`RANDOM}};
  writeStack_4_data = _RAND_60[255:0];
  _RAND_61 = {1{`RANDOM}};
  writeStack_4_mask = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  writeStack_4_validStatus = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  writeStack_4_size = _RAND_63[2:0];
  _RAND_64 = {1{`RANDOM}};
  writeStack_4_len = _RAND_64[7:0];
  _RAND_65 = {1{`RANDOM}};
  writeStack_5_wvalid = _RAND_65[0:0];
  _RAND_66 = {2{`RANDOM}};
  writeStack_5_waddr = _RAND_66[34:0];
  _RAND_67 = {1{`RANDOM}};
  writeStack_5_wstatus = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  writeStack_5_entryid = _RAND_68[4:0];
  _RAND_69 = {1{`RANDOM}};
  writeStack_5_awid = _RAND_69[13:0];
  _RAND_70 = {1{`RANDOM}};
  writeStack_5_entryFifoid = _RAND_70[4:0];
  _RAND_71 = {1{`RANDOM}};
  writeStack_5_validFifoId = _RAND_71[4:0];
  _RAND_72 = {1{`RANDOM}};
  writeStack_5_waitWFifoId = _RAND_72[4:0];
  _RAND_73 = {8{`RANDOM}};
  writeStack_5_data = _RAND_73[255:0];
  _RAND_74 = {1{`RANDOM}};
  writeStack_5_mask = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  writeStack_5_validStatus = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  writeStack_5_size = _RAND_76[2:0];
  _RAND_77 = {1{`RANDOM}};
  writeStack_5_len = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  writeStack_6_wvalid = _RAND_78[0:0];
  _RAND_79 = {2{`RANDOM}};
  writeStack_6_waddr = _RAND_79[34:0];
  _RAND_80 = {1{`RANDOM}};
  writeStack_6_wstatus = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  writeStack_6_entryid = _RAND_81[4:0];
  _RAND_82 = {1{`RANDOM}};
  writeStack_6_awid = _RAND_82[13:0];
  _RAND_83 = {1{`RANDOM}};
  writeStack_6_entryFifoid = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  writeStack_6_validFifoId = _RAND_84[4:0];
  _RAND_85 = {1{`RANDOM}};
  writeStack_6_waitWFifoId = _RAND_85[4:0];
  _RAND_86 = {8{`RANDOM}};
  writeStack_6_data = _RAND_86[255:0];
  _RAND_87 = {1{`RANDOM}};
  writeStack_6_mask = _RAND_87[31:0];
  _RAND_88 = {1{`RANDOM}};
  writeStack_6_validStatus = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  writeStack_6_size = _RAND_89[2:0];
  _RAND_90 = {1{`RANDOM}};
  writeStack_6_len = _RAND_90[7:0];
  _RAND_91 = {1{`RANDOM}};
  writeStack_7_wvalid = _RAND_91[0:0];
  _RAND_92 = {2{`RANDOM}};
  writeStack_7_waddr = _RAND_92[34:0];
  _RAND_93 = {1{`RANDOM}};
  writeStack_7_wstatus = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  writeStack_7_entryid = _RAND_94[4:0];
  _RAND_95 = {1{`RANDOM}};
  writeStack_7_awid = _RAND_95[13:0];
  _RAND_96 = {1{`RANDOM}};
  writeStack_7_entryFifoid = _RAND_96[4:0];
  _RAND_97 = {1{`RANDOM}};
  writeStack_7_validFifoId = _RAND_97[4:0];
  _RAND_98 = {1{`RANDOM}};
  writeStack_7_waitWFifoId = _RAND_98[4:0];
  _RAND_99 = {8{`RANDOM}};
  writeStack_7_data = _RAND_99[255:0];
  _RAND_100 = {1{`RANDOM}};
  writeStack_7_mask = _RAND_100[31:0];
  _RAND_101 = {1{`RANDOM}};
  writeStack_7_validStatus = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  writeStack_7_size = _RAND_102[2:0];
  _RAND_103 = {1{`RANDOM}};
  writeStack_7_len = _RAND_103[7:0];
  _RAND_104 = {1{`RANDOM}};
  writeStack_8_wvalid = _RAND_104[0:0];
  _RAND_105 = {2{`RANDOM}};
  writeStack_8_waddr = _RAND_105[34:0];
  _RAND_106 = {1{`RANDOM}};
  writeStack_8_wstatus = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  writeStack_8_entryid = _RAND_107[4:0];
  _RAND_108 = {1{`RANDOM}};
  writeStack_8_awid = _RAND_108[13:0];
  _RAND_109 = {1{`RANDOM}};
  writeStack_8_entryFifoid = _RAND_109[4:0];
  _RAND_110 = {1{`RANDOM}};
  writeStack_8_validFifoId = _RAND_110[4:0];
  _RAND_111 = {1{`RANDOM}};
  writeStack_8_waitWFifoId = _RAND_111[4:0];
  _RAND_112 = {8{`RANDOM}};
  writeStack_8_data = _RAND_112[255:0];
  _RAND_113 = {1{`RANDOM}};
  writeStack_8_mask = _RAND_113[31:0];
  _RAND_114 = {1{`RANDOM}};
  writeStack_8_validStatus = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  writeStack_8_size = _RAND_115[2:0];
  _RAND_116 = {1{`RANDOM}};
  writeStack_8_len = _RAND_116[7:0];
  _RAND_117 = {1{`RANDOM}};
  writeStack_9_wvalid = _RAND_117[0:0];
  _RAND_118 = {2{`RANDOM}};
  writeStack_9_waddr = _RAND_118[34:0];
  _RAND_119 = {1{`RANDOM}};
  writeStack_9_wstatus = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  writeStack_9_entryid = _RAND_120[4:0];
  _RAND_121 = {1{`RANDOM}};
  writeStack_9_awid = _RAND_121[13:0];
  _RAND_122 = {1{`RANDOM}};
  writeStack_9_entryFifoid = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  writeStack_9_validFifoId = _RAND_123[4:0];
  _RAND_124 = {1{`RANDOM}};
  writeStack_9_waitWFifoId = _RAND_124[4:0];
  _RAND_125 = {8{`RANDOM}};
  writeStack_9_data = _RAND_125[255:0];
  _RAND_126 = {1{`RANDOM}};
  writeStack_9_mask = _RAND_126[31:0];
  _RAND_127 = {1{`RANDOM}};
  writeStack_9_validStatus = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  writeStack_9_size = _RAND_128[2:0];
  _RAND_129 = {1{`RANDOM}};
  writeStack_9_len = _RAND_129[7:0];
  _RAND_130 = {1{`RANDOM}};
  writeStack_10_wvalid = _RAND_130[0:0];
  _RAND_131 = {2{`RANDOM}};
  writeStack_10_waddr = _RAND_131[34:0];
  _RAND_132 = {1{`RANDOM}};
  writeStack_10_wstatus = _RAND_132[1:0];
  _RAND_133 = {1{`RANDOM}};
  writeStack_10_entryid = _RAND_133[4:0];
  _RAND_134 = {1{`RANDOM}};
  writeStack_10_awid = _RAND_134[13:0];
  _RAND_135 = {1{`RANDOM}};
  writeStack_10_entryFifoid = _RAND_135[4:0];
  _RAND_136 = {1{`RANDOM}};
  writeStack_10_validFifoId = _RAND_136[4:0];
  _RAND_137 = {1{`RANDOM}};
  writeStack_10_waitWFifoId = _RAND_137[4:0];
  _RAND_138 = {8{`RANDOM}};
  writeStack_10_data = _RAND_138[255:0];
  _RAND_139 = {1{`RANDOM}};
  writeStack_10_mask = _RAND_139[31:0];
  _RAND_140 = {1{`RANDOM}};
  writeStack_10_validStatus = _RAND_140[1:0];
  _RAND_141 = {1{`RANDOM}};
  writeStack_10_size = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  writeStack_10_len = _RAND_142[7:0];
  _RAND_143 = {1{`RANDOM}};
  writeStack_11_wvalid = _RAND_143[0:0];
  _RAND_144 = {2{`RANDOM}};
  writeStack_11_waddr = _RAND_144[34:0];
  _RAND_145 = {1{`RANDOM}};
  writeStack_11_wstatus = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  writeStack_11_entryid = _RAND_146[4:0];
  _RAND_147 = {1{`RANDOM}};
  writeStack_11_awid = _RAND_147[13:0];
  _RAND_148 = {1{`RANDOM}};
  writeStack_11_entryFifoid = _RAND_148[4:0];
  _RAND_149 = {1{`RANDOM}};
  writeStack_11_validFifoId = _RAND_149[4:0];
  _RAND_150 = {1{`RANDOM}};
  writeStack_11_waitWFifoId = _RAND_150[4:0];
  _RAND_151 = {8{`RANDOM}};
  writeStack_11_data = _RAND_151[255:0];
  _RAND_152 = {1{`RANDOM}};
  writeStack_11_mask = _RAND_152[31:0];
  _RAND_153 = {1{`RANDOM}};
  writeStack_11_validStatus = _RAND_153[1:0];
  _RAND_154 = {1{`RANDOM}};
  writeStack_11_size = _RAND_154[2:0];
  _RAND_155 = {1{`RANDOM}};
  writeStack_11_len = _RAND_155[7:0];
  _RAND_156 = {1{`RANDOM}};
  writeStack_12_wvalid = _RAND_156[0:0];
  _RAND_157 = {2{`RANDOM}};
  writeStack_12_waddr = _RAND_157[34:0];
  _RAND_158 = {1{`RANDOM}};
  writeStack_12_wstatus = _RAND_158[1:0];
  _RAND_159 = {1{`RANDOM}};
  writeStack_12_entryid = _RAND_159[4:0];
  _RAND_160 = {1{`RANDOM}};
  writeStack_12_awid = _RAND_160[13:0];
  _RAND_161 = {1{`RANDOM}};
  writeStack_12_entryFifoid = _RAND_161[4:0];
  _RAND_162 = {1{`RANDOM}};
  writeStack_12_validFifoId = _RAND_162[4:0];
  _RAND_163 = {1{`RANDOM}};
  writeStack_12_waitWFifoId = _RAND_163[4:0];
  _RAND_164 = {8{`RANDOM}};
  writeStack_12_data = _RAND_164[255:0];
  _RAND_165 = {1{`RANDOM}};
  writeStack_12_mask = _RAND_165[31:0];
  _RAND_166 = {1{`RANDOM}};
  writeStack_12_validStatus = _RAND_166[1:0];
  _RAND_167 = {1{`RANDOM}};
  writeStack_12_size = _RAND_167[2:0];
  _RAND_168 = {1{`RANDOM}};
  writeStack_12_len = _RAND_168[7:0];
  _RAND_169 = {1{`RANDOM}};
  writeStack_13_wvalid = _RAND_169[0:0];
  _RAND_170 = {2{`RANDOM}};
  writeStack_13_waddr = _RAND_170[34:0];
  _RAND_171 = {1{`RANDOM}};
  writeStack_13_wstatus = _RAND_171[1:0];
  _RAND_172 = {1{`RANDOM}};
  writeStack_13_entryid = _RAND_172[4:0];
  _RAND_173 = {1{`RANDOM}};
  writeStack_13_awid = _RAND_173[13:0];
  _RAND_174 = {1{`RANDOM}};
  writeStack_13_entryFifoid = _RAND_174[4:0];
  _RAND_175 = {1{`RANDOM}};
  writeStack_13_validFifoId = _RAND_175[4:0];
  _RAND_176 = {1{`RANDOM}};
  writeStack_13_waitWFifoId = _RAND_176[4:0];
  _RAND_177 = {8{`RANDOM}};
  writeStack_13_data = _RAND_177[255:0];
  _RAND_178 = {1{`RANDOM}};
  writeStack_13_mask = _RAND_178[31:0];
  _RAND_179 = {1{`RANDOM}};
  writeStack_13_validStatus = _RAND_179[1:0];
  _RAND_180 = {1{`RANDOM}};
  writeStack_13_size = _RAND_180[2:0];
  _RAND_181 = {1{`RANDOM}};
  writeStack_13_len = _RAND_181[7:0];
  _RAND_182 = {1{`RANDOM}};
  writeStack_14_wvalid = _RAND_182[0:0];
  _RAND_183 = {2{`RANDOM}};
  writeStack_14_waddr = _RAND_183[34:0];
  _RAND_184 = {1{`RANDOM}};
  writeStack_14_wstatus = _RAND_184[1:0];
  _RAND_185 = {1{`RANDOM}};
  writeStack_14_entryid = _RAND_185[4:0];
  _RAND_186 = {1{`RANDOM}};
  writeStack_14_awid = _RAND_186[13:0];
  _RAND_187 = {1{`RANDOM}};
  writeStack_14_entryFifoid = _RAND_187[4:0];
  _RAND_188 = {1{`RANDOM}};
  writeStack_14_validFifoId = _RAND_188[4:0];
  _RAND_189 = {1{`RANDOM}};
  writeStack_14_waitWFifoId = _RAND_189[4:0];
  _RAND_190 = {8{`RANDOM}};
  writeStack_14_data = _RAND_190[255:0];
  _RAND_191 = {1{`RANDOM}};
  writeStack_14_mask = _RAND_191[31:0];
  _RAND_192 = {1{`RANDOM}};
  writeStack_14_validStatus = _RAND_192[1:0];
  _RAND_193 = {1{`RANDOM}};
  writeStack_14_size = _RAND_193[2:0];
  _RAND_194 = {1{`RANDOM}};
  writeStack_14_len = _RAND_194[7:0];
  _RAND_195 = {1{`RANDOM}};
  writeStack_15_wvalid = _RAND_195[0:0];
  _RAND_196 = {2{`RANDOM}};
  writeStack_15_waddr = _RAND_196[34:0];
  _RAND_197 = {1{`RANDOM}};
  writeStack_15_wstatus = _RAND_197[1:0];
  _RAND_198 = {1{`RANDOM}};
  writeStack_15_entryid = _RAND_198[4:0];
  _RAND_199 = {1{`RANDOM}};
  writeStack_15_awid = _RAND_199[13:0];
  _RAND_200 = {1{`RANDOM}};
  writeStack_15_entryFifoid = _RAND_200[4:0];
  _RAND_201 = {1{`RANDOM}};
  writeStack_15_validFifoId = _RAND_201[4:0];
  _RAND_202 = {1{`RANDOM}};
  writeStack_15_waitWFifoId = _RAND_202[4:0];
  _RAND_203 = {8{`RANDOM}};
  writeStack_15_data = _RAND_203[255:0];
  _RAND_204 = {1{`RANDOM}};
  writeStack_15_mask = _RAND_204[31:0];
  _RAND_205 = {1{`RANDOM}};
  writeStack_15_validStatus = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  writeStack_15_size = _RAND_206[2:0];
  _RAND_207 = {1{`RANDOM}};
  writeStack_15_len = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  writeStack_16_wvalid = _RAND_208[0:0];
  _RAND_209 = {2{`RANDOM}};
  writeStack_16_waddr = _RAND_209[34:0];
  _RAND_210 = {1{`RANDOM}};
  writeStack_16_wstatus = _RAND_210[1:0];
  _RAND_211 = {1{`RANDOM}};
  writeStack_16_entryid = _RAND_211[4:0];
  _RAND_212 = {1{`RANDOM}};
  writeStack_16_awid = _RAND_212[13:0];
  _RAND_213 = {1{`RANDOM}};
  writeStack_16_entryFifoid = _RAND_213[4:0];
  _RAND_214 = {1{`RANDOM}};
  writeStack_16_validFifoId = _RAND_214[4:0];
  _RAND_215 = {1{`RANDOM}};
  writeStack_16_waitWFifoId = _RAND_215[4:0];
  _RAND_216 = {8{`RANDOM}};
  writeStack_16_data = _RAND_216[255:0];
  _RAND_217 = {1{`RANDOM}};
  writeStack_16_mask = _RAND_217[31:0];
  _RAND_218 = {1{`RANDOM}};
  writeStack_16_validStatus = _RAND_218[1:0];
  _RAND_219 = {1{`RANDOM}};
  writeStack_16_size = _RAND_219[2:0];
  _RAND_220 = {1{`RANDOM}};
  writeStack_16_len = _RAND_220[7:0];
  _RAND_221 = {1{`RANDOM}};
  writeStack_17_wvalid = _RAND_221[0:0];
  _RAND_222 = {2{`RANDOM}};
  writeStack_17_waddr = _RAND_222[34:0];
  _RAND_223 = {1{`RANDOM}};
  writeStack_17_wstatus = _RAND_223[1:0];
  _RAND_224 = {1{`RANDOM}};
  writeStack_17_entryid = _RAND_224[4:0];
  _RAND_225 = {1{`RANDOM}};
  writeStack_17_awid = _RAND_225[13:0];
  _RAND_226 = {1{`RANDOM}};
  writeStack_17_entryFifoid = _RAND_226[4:0];
  _RAND_227 = {1{`RANDOM}};
  writeStack_17_validFifoId = _RAND_227[4:0];
  _RAND_228 = {1{`RANDOM}};
  writeStack_17_waitWFifoId = _RAND_228[4:0];
  _RAND_229 = {8{`RANDOM}};
  writeStack_17_data = _RAND_229[255:0];
  _RAND_230 = {1{`RANDOM}};
  writeStack_17_mask = _RAND_230[31:0];
  _RAND_231 = {1{`RANDOM}};
  writeStack_17_validStatus = _RAND_231[1:0];
  _RAND_232 = {1{`RANDOM}};
  writeStack_17_size = _RAND_232[2:0];
  _RAND_233 = {1{`RANDOM}};
  writeStack_17_len = _RAND_233[7:0];
  _RAND_234 = {1{`RANDOM}};
  writeStack_18_wvalid = _RAND_234[0:0];
  _RAND_235 = {2{`RANDOM}};
  writeStack_18_waddr = _RAND_235[34:0];
  _RAND_236 = {1{`RANDOM}};
  writeStack_18_wstatus = _RAND_236[1:0];
  _RAND_237 = {1{`RANDOM}};
  writeStack_18_entryid = _RAND_237[4:0];
  _RAND_238 = {1{`RANDOM}};
  writeStack_18_awid = _RAND_238[13:0];
  _RAND_239 = {1{`RANDOM}};
  writeStack_18_entryFifoid = _RAND_239[4:0];
  _RAND_240 = {1{`RANDOM}};
  writeStack_18_validFifoId = _RAND_240[4:0];
  _RAND_241 = {1{`RANDOM}};
  writeStack_18_waitWFifoId = _RAND_241[4:0];
  _RAND_242 = {8{`RANDOM}};
  writeStack_18_data = _RAND_242[255:0];
  _RAND_243 = {1{`RANDOM}};
  writeStack_18_mask = _RAND_243[31:0];
  _RAND_244 = {1{`RANDOM}};
  writeStack_18_validStatus = _RAND_244[1:0];
  _RAND_245 = {1{`RANDOM}};
  writeStack_18_size = _RAND_245[2:0];
  _RAND_246 = {1{`RANDOM}};
  writeStack_18_len = _RAND_246[7:0];
  _RAND_247 = {1{`RANDOM}};
  writeStack_19_wvalid = _RAND_247[0:0];
  _RAND_248 = {2{`RANDOM}};
  writeStack_19_waddr = _RAND_248[34:0];
  _RAND_249 = {1{`RANDOM}};
  writeStack_19_wstatus = _RAND_249[1:0];
  _RAND_250 = {1{`RANDOM}};
  writeStack_19_entryid = _RAND_250[4:0];
  _RAND_251 = {1{`RANDOM}};
  writeStack_19_awid = _RAND_251[13:0];
  _RAND_252 = {1{`RANDOM}};
  writeStack_19_entryFifoid = _RAND_252[4:0];
  _RAND_253 = {1{`RANDOM}};
  writeStack_19_validFifoId = _RAND_253[4:0];
  _RAND_254 = {1{`RANDOM}};
  writeStack_19_waitWFifoId = _RAND_254[4:0];
  _RAND_255 = {8{`RANDOM}};
  writeStack_19_data = _RAND_255[255:0];
  _RAND_256 = {1{`RANDOM}};
  writeStack_19_mask = _RAND_256[31:0];
  _RAND_257 = {1{`RANDOM}};
  writeStack_19_validStatus = _RAND_257[1:0];
  _RAND_258 = {1{`RANDOM}};
  writeStack_19_size = _RAND_258[2:0];
  _RAND_259 = {1{`RANDOM}};
  writeStack_19_len = _RAND_259[7:0];
  _RAND_260 = {1{`RANDOM}};
  writeStack_20_wvalid = _RAND_260[0:0];
  _RAND_261 = {2{`RANDOM}};
  writeStack_20_waddr = _RAND_261[34:0];
  _RAND_262 = {1{`RANDOM}};
  writeStack_20_wstatus = _RAND_262[1:0];
  _RAND_263 = {1{`RANDOM}};
  writeStack_20_entryid = _RAND_263[4:0];
  _RAND_264 = {1{`RANDOM}};
  writeStack_20_awid = _RAND_264[13:0];
  _RAND_265 = {1{`RANDOM}};
  writeStack_20_entryFifoid = _RAND_265[4:0];
  _RAND_266 = {1{`RANDOM}};
  writeStack_20_validFifoId = _RAND_266[4:0];
  _RAND_267 = {1{`RANDOM}};
  writeStack_20_waitWFifoId = _RAND_267[4:0];
  _RAND_268 = {8{`RANDOM}};
  writeStack_20_data = _RAND_268[255:0];
  _RAND_269 = {1{`RANDOM}};
  writeStack_20_mask = _RAND_269[31:0];
  _RAND_270 = {1{`RANDOM}};
  writeStack_20_validStatus = _RAND_270[1:0];
  _RAND_271 = {1{`RANDOM}};
  writeStack_20_size = _RAND_271[2:0];
  _RAND_272 = {1{`RANDOM}};
  writeStack_20_len = _RAND_272[7:0];
  _RAND_273 = {1{`RANDOM}};
  writeStack_21_wvalid = _RAND_273[0:0];
  _RAND_274 = {2{`RANDOM}};
  writeStack_21_waddr = _RAND_274[34:0];
  _RAND_275 = {1{`RANDOM}};
  writeStack_21_wstatus = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  writeStack_21_entryid = _RAND_276[4:0];
  _RAND_277 = {1{`RANDOM}};
  writeStack_21_awid = _RAND_277[13:0];
  _RAND_278 = {1{`RANDOM}};
  writeStack_21_entryFifoid = _RAND_278[4:0];
  _RAND_279 = {1{`RANDOM}};
  writeStack_21_validFifoId = _RAND_279[4:0];
  _RAND_280 = {1{`RANDOM}};
  writeStack_21_waitWFifoId = _RAND_280[4:0];
  _RAND_281 = {8{`RANDOM}};
  writeStack_21_data = _RAND_281[255:0];
  _RAND_282 = {1{`RANDOM}};
  writeStack_21_mask = _RAND_282[31:0];
  _RAND_283 = {1{`RANDOM}};
  writeStack_21_validStatus = _RAND_283[1:0];
  _RAND_284 = {1{`RANDOM}};
  writeStack_21_size = _RAND_284[2:0];
  _RAND_285 = {1{`RANDOM}};
  writeStack_21_len = _RAND_285[7:0];
  _RAND_286 = {1{`RANDOM}};
  writeStack_22_wvalid = _RAND_286[0:0];
  _RAND_287 = {2{`RANDOM}};
  writeStack_22_waddr = _RAND_287[34:0];
  _RAND_288 = {1{`RANDOM}};
  writeStack_22_wstatus = _RAND_288[1:0];
  _RAND_289 = {1{`RANDOM}};
  writeStack_22_entryid = _RAND_289[4:0];
  _RAND_290 = {1{`RANDOM}};
  writeStack_22_awid = _RAND_290[13:0];
  _RAND_291 = {1{`RANDOM}};
  writeStack_22_entryFifoid = _RAND_291[4:0];
  _RAND_292 = {1{`RANDOM}};
  writeStack_22_validFifoId = _RAND_292[4:0];
  _RAND_293 = {1{`RANDOM}};
  writeStack_22_waitWFifoId = _RAND_293[4:0];
  _RAND_294 = {8{`RANDOM}};
  writeStack_22_data = _RAND_294[255:0];
  _RAND_295 = {1{`RANDOM}};
  writeStack_22_mask = _RAND_295[31:0];
  _RAND_296 = {1{`RANDOM}};
  writeStack_22_validStatus = _RAND_296[1:0];
  _RAND_297 = {1{`RANDOM}};
  writeStack_22_size = _RAND_297[2:0];
  _RAND_298 = {1{`RANDOM}};
  writeStack_22_len = _RAND_298[7:0];
  _RAND_299 = {1{`RANDOM}};
  writeStack_23_wvalid = _RAND_299[0:0];
  _RAND_300 = {2{`RANDOM}};
  writeStack_23_waddr = _RAND_300[34:0];
  _RAND_301 = {1{`RANDOM}};
  writeStack_23_wstatus = _RAND_301[1:0];
  _RAND_302 = {1{`RANDOM}};
  writeStack_23_entryid = _RAND_302[4:0];
  _RAND_303 = {1{`RANDOM}};
  writeStack_23_awid = _RAND_303[13:0];
  _RAND_304 = {1{`RANDOM}};
  writeStack_23_entryFifoid = _RAND_304[4:0];
  _RAND_305 = {1{`RANDOM}};
  writeStack_23_validFifoId = _RAND_305[4:0];
  _RAND_306 = {1{`RANDOM}};
  writeStack_23_waitWFifoId = _RAND_306[4:0];
  _RAND_307 = {8{`RANDOM}};
  writeStack_23_data = _RAND_307[255:0];
  _RAND_308 = {1{`RANDOM}};
  writeStack_23_mask = _RAND_308[31:0];
  _RAND_309 = {1{`RANDOM}};
  writeStack_23_validStatus = _RAND_309[1:0];
  _RAND_310 = {1{`RANDOM}};
  writeStack_23_size = _RAND_310[2:0];
  _RAND_311 = {1{`RANDOM}};
  writeStack_23_len = _RAND_311[7:0];
  _RAND_312 = {1{`RANDOM}};
  writeStack_24_wvalid = _RAND_312[0:0];
  _RAND_313 = {2{`RANDOM}};
  writeStack_24_waddr = _RAND_313[34:0];
  _RAND_314 = {1{`RANDOM}};
  writeStack_24_wstatus = _RAND_314[1:0];
  _RAND_315 = {1{`RANDOM}};
  writeStack_24_entryid = _RAND_315[4:0];
  _RAND_316 = {1{`RANDOM}};
  writeStack_24_awid = _RAND_316[13:0];
  _RAND_317 = {1{`RANDOM}};
  writeStack_24_entryFifoid = _RAND_317[4:0];
  _RAND_318 = {1{`RANDOM}};
  writeStack_24_validFifoId = _RAND_318[4:0];
  _RAND_319 = {1{`RANDOM}};
  writeStack_24_waitWFifoId = _RAND_319[4:0];
  _RAND_320 = {8{`RANDOM}};
  writeStack_24_data = _RAND_320[255:0];
  _RAND_321 = {1{`RANDOM}};
  writeStack_24_mask = _RAND_321[31:0];
  _RAND_322 = {1{`RANDOM}};
  writeStack_24_validStatus = _RAND_322[1:0];
  _RAND_323 = {1{`RANDOM}};
  writeStack_24_size = _RAND_323[2:0];
  _RAND_324 = {1{`RANDOM}};
  writeStack_24_len = _RAND_324[7:0];
  _RAND_325 = {1{`RANDOM}};
  writeStack_25_wvalid = _RAND_325[0:0];
  _RAND_326 = {2{`RANDOM}};
  writeStack_25_waddr = _RAND_326[34:0];
  _RAND_327 = {1{`RANDOM}};
  writeStack_25_wstatus = _RAND_327[1:0];
  _RAND_328 = {1{`RANDOM}};
  writeStack_25_entryid = _RAND_328[4:0];
  _RAND_329 = {1{`RANDOM}};
  writeStack_25_awid = _RAND_329[13:0];
  _RAND_330 = {1{`RANDOM}};
  writeStack_25_entryFifoid = _RAND_330[4:0];
  _RAND_331 = {1{`RANDOM}};
  writeStack_25_validFifoId = _RAND_331[4:0];
  _RAND_332 = {1{`RANDOM}};
  writeStack_25_waitWFifoId = _RAND_332[4:0];
  _RAND_333 = {8{`RANDOM}};
  writeStack_25_data = _RAND_333[255:0];
  _RAND_334 = {1{`RANDOM}};
  writeStack_25_mask = _RAND_334[31:0];
  _RAND_335 = {1{`RANDOM}};
  writeStack_25_validStatus = _RAND_335[1:0];
  _RAND_336 = {1{`RANDOM}};
  writeStack_25_size = _RAND_336[2:0];
  _RAND_337 = {1{`RANDOM}};
  writeStack_25_len = _RAND_337[7:0];
  _RAND_338 = {1{`RANDOM}};
  writeStack_26_wvalid = _RAND_338[0:0];
  _RAND_339 = {2{`RANDOM}};
  writeStack_26_waddr = _RAND_339[34:0];
  _RAND_340 = {1{`RANDOM}};
  writeStack_26_wstatus = _RAND_340[1:0];
  _RAND_341 = {1{`RANDOM}};
  writeStack_26_entryid = _RAND_341[4:0];
  _RAND_342 = {1{`RANDOM}};
  writeStack_26_awid = _RAND_342[13:0];
  _RAND_343 = {1{`RANDOM}};
  writeStack_26_entryFifoid = _RAND_343[4:0];
  _RAND_344 = {1{`RANDOM}};
  writeStack_26_validFifoId = _RAND_344[4:0];
  _RAND_345 = {1{`RANDOM}};
  writeStack_26_waitWFifoId = _RAND_345[4:0];
  _RAND_346 = {8{`RANDOM}};
  writeStack_26_data = _RAND_346[255:0];
  _RAND_347 = {1{`RANDOM}};
  writeStack_26_mask = _RAND_347[31:0];
  _RAND_348 = {1{`RANDOM}};
  writeStack_26_validStatus = _RAND_348[1:0];
  _RAND_349 = {1{`RANDOM}};
  writeStack_26_size = _RAND_349[2:0];
  _RAND_350 = {1{`RANDOM}};
  writeStack_26_len = _RAND_350[7:0];
  _RAND_351 = {1{`RANDOM}};
  writeStack_27_wvalid = _RAND_351[0:0];
  _RAND_352 = {2{`RANDOM}};
  writeStack_27_waddr = _RAND_352[34:0];
  _RAND_353 = {1{`RANDOM}};
  writeStack_27_wstatus = _RAND_353[1:0];
  _RAND_354 = {1{`RANDOM}};
  writeStack_27_entryid = _RAND_354[4:0];
  _RAND_355 = {1{`RANDOM}};
  writeStack_27_awid = _RAND_355[13:0];
  _RAND_356 = {1{`RANDOM}};
  writeStack_27_entryFifoid = _RAND_356[4:0];
  _RAND_357 = {1{`RANDOM}};
  writeStack_27_validFifoId = _RAND_357[4:0];
  _RAND_358 = {1{`RANDOM}};
  writeStack_27_waitWFifoId = _RAND_358[4:0];
  _RAND_359 = {8{`RANDOM}};
  writeStack_27_data = _RAND_359[255:0];
  _RAND_360 = {1{`RANDOM}};
  writeStack_27_mask = _RAND_360[31:0];
  _RAND_361 = {1{`RANDOM}};
  writeStack_27_validStatus = _RAND_361[1:0];
  _RAND_362 = {1{`RANDOM}};
  writeStack_27_size = _RAND_362[2:0];
  _RAND_363 = {1{`RANDOM}};
  writeStack_27_len = _RAND_363[7:0];
  _RAND_364 = {1{`RANDOM}};
  writeStack_28_wvalid = _RAND_364[0:0];
  _RAND_365 = {2{`RANDOM}};
  writeStack_28_waddr = _RAND_365[34:0];
  _RAND_366 = {1{`RANDOM}};
  writeStack_28_wstatus = _RAND_366[1:0];
  _RAND_367 = {1{`RANDOM}};
  writeStack_28_entryid = _RAND_367[4:0];
  _RAND_368 = {1{`RANDOM}};
  writeStack_28_awid = _RAND_368[13:0];
  _RAND_369 = {1{`RANDOM}};
  writeStack_28_entryFifoid = _RAND_369[4:0];
  _RAND_370 = {1{`RANDOM}};
  writeStack_28_validFifoId = _RAND_370[4:0];
  _RAND_371 = {1{`RANDOM}};
  writeStack_28_waitWFifoId = _RAND_371[4:0];
  _RAND_372 = {8{`RANDOM}};
  writeStack_28_data = _RAND_372[255:0];
  _RAND_373 = {1{`RANDOM}};
  writeStack_28_mask = _RAND_373[31:0];
  _RAND_374 = {1{`RANDOM}};
  writeStack_28_validStatus = _RAND_374[1:0];
  _RAND_375 = {1{`RANDOM}};
  writeStack_28_size = _RAND_375[2:0];
  _RAND_376 = {1{`RANDOM}};
  writeStack_28_len = _RAND_376[7:0];
  _RAND_377 = {1{`RANDOM}};
  writeStack_29_wvalid = _RAND_377[0:0];
  _RAND_378 = {2{`RANDOM}};
  writeStack_29_waddr = _RAND_378[34:0];
  _RAND_379 = {1{`RANDOM}};
  writeStack_29_wstatus = _RAND_379[1:0];
  _RAND_380 = {1{`RANDOM}};
  writeStack_29_entryid = _RAND_380[4:0];
  _RAND_381 = {1{`RANDOM}};
  writeStack_29_awid = _RAND_381[13:0];
  _RAND_382 = {1{`RANDOM}};
  writeStack_29_entryFifoid = _RAND_382[4:0];
  _RAND_383 = {1{`RANDOM}};
  writeStack_29_validFifoId = _RAND_383[4:0];
  _RAND_384 = {1{`RANDOM}};
  writeStack_29_waitWFifoId = _RAND_384[4:0];
  _RAND_385 = {8{`RANDOM}};
  writeStack_29_data = _RAND_385[255:0];
  _RAND_386 = {1{`RANDOM}};
  writeStack_29_mask = _RAND_386[31:0];
  _RAND_387 = {1{`RANDOM}};
  writeStack_29_validStatus = _RAND_387[1:0];
  _RAND_388 = {1{`RANDOM}};
  writeStack_29_size = _RAND_388[2:0];
  _RAND_389 = {1{`RANDOM}};
  writeStack_29_len = _RAND_389[7:0];
  _RAND_390 = {1{`RANDOM}};
  writeStack_30_wvalid = _RAND_390[0:0];
  _RAND_391 = {2{`RANDOM}};
  writeStack_30_waddr = _RAND_391[34:0];
  _RAND_392 = {1{`RANDOM}};
  writeStack_30_wstatus = _RAND_392[1:0];
  _RAND_393 = {1{`RANDOM}};
  writeStack_30_entryid = _RAND_393[4:0];
  _RAND_394 = {1{`RANDOM}};
  writeStack_30_awid = _RAND_394[13:0];
  _RAND_395 = {1{`RANDOM}};
  writeStack_30_entryFifoid = _RAND_395[4:0];
  _RAND_396 = {1{`RANDOM}};
  writeStack_30_validFifoId = _RAND_396[4:0];
  _RAND_397 = {1{`RANDOM}};
  writeStack_30_waitWFifoId = _RAND_397[4:0];
  _RAND_398 = {8{`RANDOM}};
  writeStack_30_data = _RAND_398[255:0];
  _RAND_399 = {1{`RANDOM}};
  writeStack_30_mask = _RAND_399[31:0];
  _RAND_400 = {1{`RANDOM}};
  writeStack_30_validStatus = _RAND_400[1:0];
  _RAND_401 = {1{`RANDOM}};
  writeStack_30_size = _RAND_401[2:0];
  _RAND_402 = {1{`RANDOM}};
  writeStack_30_len = _RAND_402[7:0];
  _RAND_403 = {1{`RANDOM}};
  writeStack_31_wvalid = _RAND_403[0:0];
  _RAND_404 = {2{`RANDOM}};
  writeStack_31_waddr = _RAND_404[34:0];
  _RAND_405 = {1{`RANDOM}};
  writeStack_31_wstatus = _RAND_405[1:0];
  _RAND_406 = {1{`RANDOM}};
  writeStack_31_entryid = _RAND_406[4:0];
  _RAND_407 = {1{`RANDOM}};
  writeStack_31_awid = _RAND_407[13:0];
  _RAND_408 = {1{`RANDOM}};
  writeStack_31_entryFifoid = _RAND_408[4:0];
  _RAND_409 = {1{`RANDOM}};
  writeStack_31_validFifoId = _RAND_409[4:0];
  _RAND_410 = {1{`RANDOM}};
  writeStack_31_waitWFifoId = _RAND_410[4:0];
  _RAND_411 = {8{`RANDOM}};
  writeStack_31_data = _RAND_411[255:0];
  _RAND_412 = {1{`RANDOM}};
  writeStack_31_mask = _RAND_412[31:0];
  _RAND_413 = {1{`RANDOM}};
  writeStack_31_validStatus = _RAND_413[1:0];
  _RAND_414 = {1{`RANDOM}};
  writeStack_31_size = _RAND_414[2:0];
  _RAND_415 = {1{`RANDOM}};
  writeStack_31_len = _RAND_415[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
