module Arbiter(
  input          io_in_0_valid,
  input  [34:0]  io_in_0_bits_raddress,
  input  [4:0]   io_in_0_bits_entryid,
  input  [13:0]  io_in_0_bits_arid,
  input  [255:0] io_in_0_bits_ardata,
  input  [3:0]   io_in_0_bits_respStatus,
  input  [7:0]   io_in_0_bits_rsize,
  input          io_in_1_valid,
  input  [34:0]  io_in_1_bits_raddress,
  input  [4:0]   io_in_1_bits_entryid,
  input  [13:0]  io_in_1_bits_arid,
  input  [255:0] io_in_1_bits_ardata,
  input  [3:0]   io_in_1_bits_respStatus,
  input  [7:0]   io_in_1_bits_rsize,
  input          io_in_2_valid,
  input  [34:0]  io_in_2_bits_raddress,
  input  [4:0]   io_in_2_bits_entryid,
  input  [13:0]  io_in_2_bits_arid,
  input  [255:0] io_in_2_bits_ardata,
  input  [3:0]   io_in_2_bits_respStatus,
  input  [7:0]   io_in_2_bits_rsize,
  input          io_in_3_valid,
  input  [34:0]  io_in_3_bits_raddress,
  input  [4:0]   io_in_3_bits_entryid,
  input  [13:0]  io_in_3_bits_arid,
  input  [255:0] io_in_3_bits_ardata,
  input  [3:0]   io_in_3_bits_respStatus,
  input  [7:0]   io_in_3_bits_rsize,
  input          io_in_4_valid,
  input  [34:0]  io_in_4_bits_raddress,
  input  [4:0]   io_in_4_bits_entryid,
  input  [13:0]  io_in_4_bits_arid,
  input  [255:0] io_in_4_bits_ardata,
  input  [3:0]   io_in_4_bits_respStatus,
  input  [7:0]   io_in_4_bits_rsize,
  input          io_in_5_valid,
  input  [34:0]  io_in_5_bits_raddress,
  input  [4:0]   io_in_5_bits_entryid,
  input  [13:0]  io_in_5_bits_arid,
  input  [255:0] io_in_5_bits_ardata,
  input  [3:0]   io_in_5_bits_respStatus,
  input  [7:0]   io_in_5_bits_rsize,
  input          io_in_6_valid,
  input  [34:0]  io_in_6_bits_raddress,
  input  [4:0]   io_in_6_bits_entryid,
  input  [13:0]  io_in_6_bits_arid,
  input  [255:0] io_in_6_bits_ardata,
  input  [3:0]   io_in_6_bits_respStatus,
  input  [7:0]   io_in_6_bits_rsize,
  input          io_in_7_valid,
  input  [34:0]  io_in_7_bits_raddress,
  input  [4:0]   io_in_7_bits_entryid,
  input  [13:0]  io_in_7_bits_arid,
  input  [255:0] io_in_7_bits_ardata,
  input  [3:0]   io_in_7_bits_respStatus,
  input  [7:0]   io_in_7_bits_rsize,
  input          io_in_8_valid,
  input  [34:0]  io_in_8_bits_raddress,
  input  [4:0]   io_in_8_bits_entryid,
  input  [13:0]  io_in_8_bits_arid,
  input  [255:0] io_in_8_bits_ardata,
  input  [3:0]   io_in_8_bits_respStatus,
  input  [7:0]   io_in_8_bits_rsize,
  input          io_in_9_valid,
  input  [34:0]  io_in_9_bits_raddress,
  input  [4:0]   io_in_9_bits_entryid,
  input  [13:0]  io_in_9_bits_arid,
  input  [255:0] io_in_9_bits_ardata,
  input  [3:0]   io_in_9_bits_respStatus,
  input  [7:0]   io_in_9_bits_rsize,
  input          io_in_10_valid,
  input  [34:0]  io_in_10_bits_raddress,
  input  [4:0]   io_in_10_bits_entryid,
  input  [13:0]  io_in_10_bits_arid,
  input  [255:0] io_in_10_bits_ardata,
  input  [3:0]   io_in_10_bits_respStatus,
  input  [7:0]   io_in_10_bits_rsize,
  input          io_in_11_valid,
  input  [34:0]  io_in_11_bits_raddress,
  input  [4:0]   io_in_11_bits_entryid,
  input  [13:0]  io_in_11_bits_arid,
  input  [255:0] io_in_11_bits_ardata,
  input  [3:0]   io_in_11_bits_respStatus,
  input  [7:0]   io_in_11_bits_rsize,
  input          io_in_12_valid,
  input  [34:0]  io_in_12_bits_raddress,
  input  [4:0]   io_in_12_bits_entryid,
  input  [13:0]  io_in_12_bits_arid,
  input  [255:0] io_in_12_bits_ardata,
  input  [3:0]   io_in_12_bits_respStatus,
  input  [7:0]   io_in_12_bits_rsize,
  input          io_in_13_valid,
  input  [34:0]  io_in_13_bits_raddress,
  input  [4:0]   io_in_13_bits_entryid,
  input  [13:0]  io_in_13_bits_arid,
  input  [255:0] io_in_13_bits_ardata,
  input  [3:0]   io_in_13_bits_respStatus,
  input  [7:0]   io_in_13_bits_rsize,
  input          io_in_14_valid,
  input  [34:0]  io_in_14_bits_raddress,
  input  [4:0]   io_in_14_bits_entryid,
  input  [13:0]  io_in_14_bits_arid,
  input  [255:0] io_in_14_bits_ardata,
  input  [3:0]   io_in_14_bits_respStatus,
  input  [7:0]   io_in_14_bits_rsize,
  input          io_in_15_valid,
  input  [34:0]  io_in_15_bits_raddress,
  input  [4:0]   io_in_15_bits_entryid,
  input  [13:0]  io_in_15_bits_arid,
  input  [255:0] io_in_15_bits_ardata,
  input  [3:0]   io_in_15_bits_respStatus,
  input  [7:0]   io_in_15_bits_rsize,
  input          io_in_16_valid,
  input  [34:0]  io_in_16_bits_raddress,
  input  [4:0]   io_in_16_bits_entryid,
  input  [13:0]  io_in_16_bits_arid,
  input  [255:0] io_in_16_bits_ardata,
  input  [3:0]   io_in_16_bits_respStatus,
  input  [7:0]   io_in_16_bits_rsize,
  input          io_in_17_valid,
  input  [34:0]  io_in_17_bits_raddress,
  input  [4:0]   io_in_17_bits_entryid,
  input  [13:0]  io_in_17_bits_arid,
  input  [255:0] io_in_17_bits_ardata,
  input  [3:0]   io_in_17_bits_respStatus,
  input  [7:0]   io_in_17_bits_rsize,
  input          io_in_18_valid,
  input  [34:0]  io_in_18_bits_raddress,
  input  [4:0]   io_in_18_bits_entryid,
  input  [13:0]  io_in_18_bits_arid,
  input  [255:0] io_in_18_bits_ardata,
  input  [3:0]   io_in_18_bits_respStatus,
  input  [7:0]   io_in_18_bits_rsize,
  input          io_in_19_valid,
  input  [34:0]  io_in_19_bits_raddress,
  input  [4:0]   io_in_19_bits_entryid,
  input  [13:0]  io_in_19_bits_arid,
  input  [255:0] io_in_19_bits_ardata,
  input  [3:0]   io_in_19_bits_respStatus,
  input  [7:0]   io_in_19_bits_rsize,
  input          io_in_20_valid,
  input  [34:0]  io_in_20_bits_raddress,
  input  [4:0]   io_in_20_bits_entryid,
  input  [13:0]  io_in_20_bits_arid,
  input  [255:0] io_in_20_bits_ardata,
  input  [3:0]   io_in_20_bits_respStatus,
  input  [7:0]   io_in_20_bits_rsize,
  input          io_in_21_valid,
  input  [34:0]  io_in_21_bits_raddress,
  input  [4:0]   io_in_21_bits_entryid,
  input  [13:0]  io_in_21_bits_arid,
  input  [255:0] io_in_21_bits_ardata,
  input  [3:0]   io_in_21_bits_respStatus,
  input  [7:0]   io_in_21_bits_rsize,
  input          io_in_22_valid,
  input  [34:0]  io_in_22_bits_raddress,
  input  [4:0]   io_in_22_bits_entryid,
  input  [13:0]  io_in_22_bits_arid,
  input  [255:0] io_in_22_bits_ardata,
  input  [3:0]   io_in_22_bits_respStatus,
  input  [7:0]   io_in_22_bits_rsize,
  input          io_in_23_valid,
  input  [34:0]  io_in_23_bits_raddress,
  input  [4:0]   io_in_23_bits_entryid,
  input  [13:0]  io_in_23_bits_arid,
  input  [255:0] io_in_23_bits_ardata,
  input  [3:0]   io_in_23_bits_respStatus,
  input  [7:0]   io_in_23_bits_rsize,
  input          io_in_24_valid,
  input  [34:0]  io_in_24_bits_raddress,
  input  [4:0]   io_in_24_bits_entryid,
  input  [13:0]  io_in_24_bits_arid,
  input  [255:0] io_in_24_bits_ardata,
  input  [3:0]   io_in_24_bits_respStatus,
  input  [7:0]   io_in_24_bits_rsize,
  input          io_in_25_valid,
  input  [34:0]  io_in_25_bits_raddress,
  input  [4:0]   io_in_25_bits_entryid,
  input  [13:0]  io_in_25_bits_arid,
  input  [255:0] io_in_25_bits_ardata,
  input  [3:0]   io_in_25_bits_respStatus,
  input  [7:0]   io_in_25_bits_rsize,
  input          io_in_26_valid,
  input  [34:0]  io_in_26_bits_raddress,
  input  [4:0]   io_in_26_bits_entryid,
  input  [13:0]  io_in_26_bits_arid,
  input  [255:0] io_in_26_bits_ardata,
  input  [3:0]   io_in_26_bits_respStatus,
  input  [7:0]   io_in_26_bits_rsize,
  input          io_in_27_valid,
  input  [34:0]  io_in_27_bits_raddress,
  input  [4:0]   io_in_27_bits_entryid,
  input  [13:0]  io_in_27_bits_arid,
  input  [255:0] io_in_27_bits_ardata,
  input  [3:0]   io_in_27_bits_respStatus,
  input  [7:0]   io_in_27_bits_rsize,
  input          io_in_28_valid,
  input  [34:0]  io_in_28_bits_raddress,
  input  [4:0]   io_in_28_bits_entryid,
  input  [13:0]  io_in_28_bits_arid,
  input  [255:0] io_in_28_bits_ardata,
  input  [3:0]   io_in_28_bits_respStatus,
  input  [7:0]   io_in_28_bits_rsize,
  input          io_in_29_valid,
  input  [34:0]  io_in_29_bits_raddress,
  input  [4:0]   io_in_29_bits_entryid,
  input  [13:0]  io_in_29_bits_arid,
  input  [255:0] io_in_29_bits_ardata,
  input  [3:0]   io_in_29_bits_respStatus,
  input  [7:0]   io_in_29_bits_rsize,
  input          io_in_30_valid,
  input  [34:0]  io_in_30_bits_raddress,
  input  [4:0]   io_in_30_bits_entryid,
  input  [13:0]  io_in_30_bits_arid,
  input  [255:0] io_in_30_bits_ardata,
  input  [3:0]   io_in_30_bits_respStatus,
  input  [7:0]   io_in_30_bits_rsize,
  input          io_in_31_valid,
  input  [34:0]  io_in_31_bits_raddress,
  input  [4:0]   io_in_31_bits_entryid,
  input  [13:0]  io_in_31_bits_arid,
  input  [255:0] io_in_31_bits_ardata,
  input  [3:0]   io_in_31_bits_respStatus,
  input  [7:0]   io_in_31_bits_rsize,
  output         io_out_valid,
  output [34:0]  io_out_bits_raddress,
  output [4:0]   io_out_bits_entryid,
  output [13:0]  io_out_bits_arid,
  output [255:0] io_out_bits_ardata,
  output [3:0]   io_out_bits_respStatus,
  output [7:0]   io_out_bits_rsize,
  output [4:0]   io_chosen
);
  wire [4:0] _GEN_0 = io_in_30_valid ? 5'h1e : 5'h1f; // @[Arbiter.scala 138:13 141:26 142:17]
  wire [7:0] _GEN_6 = io_in_30_valid ? io_in_30_bits_rsize : io_in_31_bits_rsize; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [3:0] _GEN_7 = io_in_30_valid ? io_in_30_bits_respStatus : io_in_31_bits_respStatus; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [255:0] _GEN_9 = io_in_30_valid ? io_in_30_bits_ardata : io_in_31_bits_ardata; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [13:0] _GEN_10 = io_in_30_valid ? io_in_30_bits_arid : io_in_31_bits_arid; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [4:0] _GEN_11 = io_in_30_valid ? io_in_30_bits_entryid : io_in_31_bits_entryid; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [34:0] _GEN_12 = io_in_30_valid ? io_in_30_bits_raddress : io_in_31_bits_raddress; // @[Arbiter.scala 139:15 141:26 143:19]
  wire [4:0] _GEN_15 = io_in_29_valid ? 5'h1d : _GEN_0; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_21 = io_in_29_valid ? io_in_29_bits_rsize : _GEN_6; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_22 = io_in_29_valid ? io_in_29_bits_respStatus : _GEN_7; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_24 = io_in_29_valid ? io_in_29_bits_ardata : _GEN_9; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_25 = io_in_29_valid ? io_in_29_bits_arid : _GEN_10; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_26 = io_in_29_valid ? io_in_29_bits_entryid : _GEN_11; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_27 = io_in_29_valid ? io_in_29_bits_raddress : _GEN_12; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_30 = io_in_28_valid ? 5'h1c : _GEN_15; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_36 = io_in_28_valid ? io_in_28_bits_rsize : _GEN_21; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_37 = io_in_28_valid ? io_in_28_bits_respStatus : _GEN_22; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_39 = io_in_28_valid ? io_in_28_bits_ardata : _GEN_24; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_40 = io_in_28_valid ? io_in_28_bits_arid : _GEN_25; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_41 = io_in_28_valid ? io_in_28_bits_entryid : _GEN_26; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_42 = io_in_28_valid ? io_in_28_bits_raddress : _GEN_27; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_45 = io_in_27_valid ? 5'h1b : _GEN_30; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_51 = io_in_27_valid ? io_in_27_bits_rsize : _GEN_36; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_52 = io_in_27_valid ? io_in_27_bits_respStatus : _GEN_37; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_54 = io_in_27_valid ? io_in_27_bits_ardata : _GEN_39; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_55 = io_in_27_valid ? io_in_27_bits_arid : _GEN_40; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_56 = io_in_27_valid ? io_in_27_bits_entryid : _GEN_41; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_57 = io_in_27_valid ? io_in_27_bits_raddress : _GEN_42; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_60 = io_in_26_valid ? 5'h1a : _GEN_45; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_66 = io_in_26_valid ? io_in_26_bits_rsize : _GEN_51; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_67 = io_in_26_valid ? io_in_26_bits_respStatus : _GEN_52; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_69 = io_in_26_valid ? io_in_26_bits_ardata : _GEN_54; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_70 = io_in_26_valid ? io_in_26_bits_arid : _GEN_55; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_71 = io_in_26_valid ? io_in_26_bits_entryid : _GEN_56; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_72 = io_in_26_valid ? io_in_26_bits_raddress : _GEN_57; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_75 = io_in_25_valid ? 5'h19 : _GEN_60; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_81 = io_in_25_valid ? io_in_25_bits_rsize : _GEN_66; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_82 = io_in_25_valid ? io_in_25_bits_respStatus : _GEN_67; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_84 = io_in_25_valid ? io_in_25_bits_ardata : _GEN_69; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_85 = io_in_25_valid ? io_in_25_bits_arid : _GEN_70; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_86 = io_in_25_valid ? io_in_25_bits_entryid : _GEN_71; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_87 = io_in_25_valid ? io_in_25_bits_raddress : _GEN_72; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_90 = io_in_24_valid ? 5'h18 : _GEN_75; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_96 = io_in_24_valid ? io_in_24_bits_rsize : _GEN_81; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_97 = io_in_24_valid ? io_in_24_bits_respStatus : _GEN_82; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_99 = io_in_24_valid ? io_in_24_bits_ardata : _GEN_84; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_100 = io_in_24_valid ? io_in_24_bits_arid : _GEN_85; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_101 = io_in_24_valid ? io_in_24_bits_entryid : _GEN_86; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_102 = io_in_24_valid ? io_in_24_bits_raddress : _GEN_87; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_105 = io_in_23_valid ? 5'h17 : _GEN_90; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_111 = io_in_23_valid ? io_in_23_bits_rsize : _GEN_96; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_112 = io_in_23_valid ? io_in_23_bits_respStatus : _GEN_97; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_114 = io_in_23_valid ? io_in_23_bits_ardata : _GEN_99; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_115 = io_in_23_valid ? io_in_23_bits_arid : _GEN_100; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_116 = io_in_23_valid ? io_in_23_bits_entryid : _GEN_101; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_117 = io_in_23_valid ? io_in_23_bits_raddress : _GEN_102; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_120 = io_in_22_valid ? 5'h16 : _GEN_105; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_126 = io_in_22_valid ? io_in_22_bits_rsize : _GEN_111; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_127 = io_in_22_valid ? io_in_22_bits_respStatus : _GEN_112; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_129 = io_in_22_valid ? io_in_22_bits_ardata : _GEN_114; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_130 = io_in_22_valid ? io_in_22_bits_arid : _GEN_115; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_131 = io_in_22_valid ? io_in_22_bits_entryid : _GEN_116; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_132 = io_in_22_valid ? io_in_22_bits_raddress : _GEN_117; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_135 = io_in_21_valid ? 5'h15 : _GEN_120; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_141 = io_in_21_valid ? io_in_21_bits_rsize : _GEN_126; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_142 = io_in_21_valid ? io_in_21_bits_respStatus : _GEN_127; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_144 = io_in_21_valid ? io_in_21_bits_ardata : _GEN_129; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_145 = io_in_21_valid ? io_in_21_bits_arid : _GEN_130; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_146 = io_in_21_valid ? io_in_21_bits_entryid : _GEN_131; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_147 = io_in_21_valid ? io_in_21_bits_raddress : _GEN_132; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_150 = io_in_20_valid ? 5'h14 : _GEN_135; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_156 = io_in_20_valid ? io_in_20_bits_rsize : _GEN_141; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_157 = io_in_20_valid ? io_in_20_bits_respStatus : _GEN_142; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_159 = io_in_20_valid ? io_in_20_bits_ardata : _GEN_144; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_160 = io_in_20_valid ? io_in_20_bits_arid : _GEN_145; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_161 = io_in_20_valid ? io_in_20_bits_entryid : _GEN_146; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_162 = io_in_20_valid ? io_in_20_bits_raddress : _GEN_147; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_165 = io_in_19_valid ? 5'h13 : _GEN_150; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_171 = io_in_19_valid ? io_in_19_bits_rsize : _GEN_156; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_172 = io_in_19_valid ? io_in_19_bits_respStatus : _GEN_157; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_174 = io_in_19_valid ? io_in_19_bits_ardata : _GEN_159; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_175 = io_in_19_valid ? io_in_19_bits_arid : _GEN_160; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_176 = io_in_19_valid ? io_in_19_bits_entryid : _GEN_161; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_177 = io_in_19_valid ? io_in_19_bits_raddress : _GEN_162; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_180 = io_in_18_valid ? 5'h12 : _GEN_165; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_186 = io_in_18_valid ? io_in_18_bits_rsize : _GEN_171; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_187 = io_in_18_valid ? io_in_18_bits_respStatus : _GEN_172; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_189 = io_in_18_valid ? io_in_18_bits_ardata : _GEN_174; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_190 = io_in_18_valid ? io_in_18_bits_arid : _GEN_175; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_191 = io_in_18_valid ? io_in_18_bits_entryid : _GEN_176; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_192 = io_in_18_valid ? io_in_18_bits_raddress : _GEN_177; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_195 = io_in_17_valid ? 5'h11 : _GEN_180; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_201 = io_in_17_valid ? io_in_17_bits_rsize : _GEN_186; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_202 = io_in_17_valid ? io_in_17_bits_respStatus : _GEN_187; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_204 = io_in_17_valid ? io_in_17_bits_ardata : _GEN_189; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_205 = io_in_17_valid ? io_in_17_bits_arid : _GEN_190; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_206 = io_in_17_valid ? io_in_17_bits_entryid : _GEN_191; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_207 = io_in_17_valid ? io_in_17_bits_raddress : _GEN_192; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_210 = io_in_16_valid ? 5'h10 : _GEN_195; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_216 = io_in_16_valid ? io_in_16_bits_rsize : _GEN_201; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_217 = io_in_16_valid ? io_in_16_bits_respStatus : _GEN_202; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_219 = io_in_16_valid ? io_in_16_bits_ardata : _GEN_204; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_220 = io_in_16_valid ? io_in_16_bits_arid : _GEN_205; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_221 = io_in_16_valid ? io_in_16_bits_entryid : _GEN_206; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_222 = io_in_16_valid ? io_in_16_bits_raddress : _GEN_207; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_225 = io_in_15_valid ? 5'hf : _GEN_210; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_231 = io_in_15_valid ? io_in_15_bits_rsize : _GEN_216; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_232 = io_in_15_valid ? io_in_15_bits_respStatus : _GEN_217; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_234 = io_in_15_valid ? io_in_15_bits_ardata : _GEN_219; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_235 = io_in_15_valid ? io_in_15_bits_arid : _GEN_220; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_236 = io_in_15_valid ? io_in_15_bits_entryid : _GEN_221; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_237 = io_in_15_valid ? io_in_15_bits_raddress : _GEN_222; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_240 = io_in_14_valid ? 5'he : _GEN_225; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_246 = io_in_14_valid ? io_in_14_bits_rsize : _GEN_231; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_247 = io_in_14_valid ? io_in_14_bits_respStatus : _GEN_232; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_249 = io_in_14_valid ? io_in_14_bits_ardata : _GEN_234; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_250 = io_in_14_valid ? io_in_14_bits_arid : _GEN_235; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_251 = io_in_14_valid ? io_in_14_bits_entryid : _GEN_236; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_252 = io_in_14_valid ? io_in_14_bits_raddress : _GEN_237; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_255 = io_in_13_valid ? 5'hd : _GEN_240; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_261 = io_in_13_valid ? io_in_13_bits_rsize : _GEN_246; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_262 = io_in_13_valid ? io_in_13_bits_respStatus : _GEN_247; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_264 = io_in_13_valid ? io_in_13_bits_ardata : _GEN_249; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_265 = io_in_13_valid ? io_in_13_bits_arid : _GEN_250; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_266 = io_in_13_valid ? io_in_13_bits_entryid : _GEN_251; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_267 = io_in_13_valid ? io_in_13_bits_raddress : _GEN_252; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_270 = io_in_12_valid ? 5'hc : _GEN_255; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_276 = io_in_12_valid ? io_in_12_bits_rsize : _GEN_261; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_277 = io_in_12_valid ? io_in_12_bits_respStatus : _GEN_262; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_279 = io_in_12_valid ? io_in_12_bits_ardata : _GEN_264; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_280 = io_in_12_valid ? io_in_12_bits_arid : _GEN_265; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_281 = io_in_12_valid ? io_in_12_bits_entryid : _GEN_266; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_282 = io_in_12_valid ? io_in_12_bits_raddress : _GEN_267; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_285 = io_in_11_valid ? 5'hb : _GEN_270; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_291 = io_in_11_valid ? io_in_11_bits_rsize : _GEN_276; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_292 = io_in_11_valid ? io_in_11_bits_respStatus : _GEN_277; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_294 = io_in_11_valid ? io_in_11_bits_ardata : _GEN_279; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_295 = io_in_11_valid ? io_in_11_bits_arid : _GEN_280; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_296 = io_in_11_valid ? io_in_11_bits_entryid : _GEN_281; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_297 = io_in_11_valid ? io_in_11_bits_raddress : _GEN_282; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_300 = io_in_10_valid ? 5'ha : _GEN_285; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_306 = io_in_10_valid ? io_in_10_bits_rsize : _GEN_291; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_307 = io_in_10_valid ? io_in_10_bits_respStatus : _GEN_292; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_309 = io_in_10_valid ? io_in_10_bits_ardata : _GEN_294; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_310 = io_in_10_valid ? io_in_10_bits_arid : _GEN_295; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_311 = io_in_10_valid ? io_in_10_bits_entryid : _GEN_296; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_312 = io_in_10_valid ? io_in_10_bits_raddress : _GEN_297; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_315 = io_in_9_valid ? 5'h9 : _GEN_300; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_321 = io_in_9_valid ? io_in_9_bits_rsize : _GEN_306; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_322 = io_in_9_valid ? io_in_9_bits_respStatus : _GEN_307; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_324 = io_in_9_valid ? io_in_9_bits_ardata : _GEN_309; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_325 = io_in_9_valid ? io_in_9_bits_arid : _GEN_310; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_326 = io_in_9_valid ? io_in_9_bits_entryid : _GEN_311; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_327 = io_in_9_valid ? io_in_9_bits_raddress : _GEN_312; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_330 = io_in_8_valid ? 5'h8 : _GEN_315; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_336 = io_in_8_valid ? io_in_8_bits_rsize : _GEN_321; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_337 = io_in_8_valid ? io_in_8_bits_respStatus : _GEN_322; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_339 = io_in_8_valid ? io_in_8_bits_ardata : _GEN_324; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_340 = io_in_8_valid ? io_in_8_bits_arid : _GEN_325; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_341 = io_in_8_valid ? io_in_8_bits_entryid : _GEN_326; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_342 = io_in_8_valid ? io_in_8_bits_raddress : _GEN_327; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_345 = io_in_7_valid ? 5'h7 : _GEN_330; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_351 = io_in_7_valid ? io_in_7_bits_rsize : _GEN_336; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_352 = io_in_7_valid ? io_in_7_bits_respStatus : _GEN_337; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_354 = io_in_7_valid ? io_in_7_bits_ardata : _GEN_339; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_355 = io_in_7_valid ? io_in_7_bits_arid : _GEN_340; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_356 = io_in_7_valid ? io_in_7_bits_entryid : _GEN_341; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_357 = io_in_7_valid ? io_in_7_bits_raddress : _GEN_342; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_360 = io_in_6_valid ? 5'h6 : _GEN_345; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_366 = io_in_6_valid ? io_in_6_bits_rsize : _GEN_351; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_367 = io_in_6_valid ? io_in_6_bits_respStatus : _GEN_352; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_369 = io_in_6_valid ? io_in_6_bits_ardata : _GEN_354; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_370 = io_in_6_valid ? io_in_6_bits_arid : _GEN_355; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_371 = io_in_6_valid ? io_in_6_bits_entryid : _GEN_356; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_372 = io_in_6_valid ? io_in_6_bits_raddress : _GEN_357; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_375 = io_in_5_valid ? 5'h5 : _GEN_360; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_381 = io_in_5_valid ? io_in_5_bits_rsize : _GEN_366; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_382 = io_in_5_valid ? io_in_5_bits_respStatus : _GEN_367; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_384 = io_in_5_valid ? io_in_5_bits_ardata : _GEN_369; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_385 = io_in_5_valid ? io_in_5_bits_arid : _GEN_370; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_386 = io_in_5_valid ? io_in_5_bits_entryid : _GEN_371; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_387 = io_in_5_valid ? io_in_5_bits_raddress : _GEN_372; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_390 = io_in_4_valid ? 5'h4 : _GEN_375; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_396 = io_in_4_valid ? io_in_4_bits_rsize : _GEN_381; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_397 = io_in_4_valid ? io_in_4_bits_respStatus : _GEN_382; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_399 = io_in_4_valid ? io_in_4_bits_ardata : _GEN_384; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_400 = io_in_4_valid ? io_in_4_bits_arid : _GEN_385; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_401 = io_in_4_valid ? io_in_4_bits_entryid : _GEN_386; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_402 = io_in_4_valid ? io_in_4_bits_raddress : _GEN_387; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_405 = io_in_3_valid ? 5'h3 : _GEN_390; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_411 = io_in_3_valid ? io_in_3_bits_rsize : _GEN_396; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_412 = io_in_3_valid ? io_in_3_bits_respStatus : _GEN_397; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_414 = io_in_3_valid ? io_in_3_bits_ardata : _GEN_399; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_415 = io_in_3_valid ? io_in_3_bits_arid : _GEN_400; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_416 = io_in_3_valid ? io_in_3_bits_entryid : _GEN_401; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_417 = io_in_3_valid ? io_in_3_bits_raddress : _GEN_402; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_420 = io_in_2_valid ? 5'h2 : _GEN_405; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_426 = io_in_2_valid ? io_in_2_bits_rsize : _GEN_411; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_427 = io_in_2_valid ? io_in_2_bits_respStatus : _GEN_412; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_429 = io_in_2_valid ? io_in_2_bits_ardata : _GEN_414; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_430 = io_in_2_valid ? io_in_2_bits_arid : _GEN_415; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_431 = io_in_2_valid ? io_in_2_bits_entryid : _GEN_416; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_432 = io_in_2_valid ? io_in_2_bits_raddress : _GEN_417; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_435 = io_in_1_valid ? 5'h1 : _GEN_420; // @[Arbiter.scala 141:26 142:17]
  wire [7:0] _GEN_441 = io_in_1_valid ? io_in_1_bits_rsize : _GEN_426; // @[Arbiter.scala 141:26 143:19]
  wire [3:0] _GEN_442 = io_in_1_valid ? io_in_1_bits_respStatus : _GEN_427; // @[Arbiter.scala 141:26 143:19]
  wire [255:0] _GEN_444 = io_in_1_valid ? io_in_1_bits_ardata : _GEN_429; // @[Arbiter.scala 141:26 143:19]
  wire [13:0] _GEN_445 = io_in_1_valid ? io_in_1_bits_arid : _GEN_430; // @[Arbiter.scala 141:26 143:19]
  wire [4:0] _GEN_446 = io_in_1_valid ? io_in_1_bits_entryid : _GEN_431; // @[Arbiter.scala 141:26 143:19]
  wire [34:0] _GEN_447 = io_in_1_valid ? io_in_1_bits_raddress : _GEN_432; // @[Arbiter.scala 141:26 143:19]
  wire  _grant_T_29 = io_in_0_valid | io_in_1_valid | io_in_2_valid | io_in_3_valid | io_in_4_valid | io_in_5_valid |
    io_in_6_valid | io_in_7_valid | io_in_8_valid | io_in_9_valid | io_in_10_valid | io_in_11_valid | io_in_12_valid |
    io_in_13_valid | io_in_14_valid | io_in_15_valid | io_in_16_valid | io_in_17_valid | io_in_18_valid | io_in_19_valid
     | io_in_20_valid | io_in_21_valid | io_in_22_valid | io_in_23_valid | io_in_24_valid | io_in_25_valid |
    io_in_26_valid | io_in_27_valid | io_in_28_valid | io_in_29_valid | io_in_30_valid; // @[Arbiter.scala 46:68]
  wire  grant_31 = ~_grant_T_29; // @[Arbiter.scala 46:78]
  assign io_out_valid = ~grant_31 | io_in_31_valid; // @[Arbiter.scala 150:31]
  assign io_out_bits_raddress = io_in_0_valid ? io_in_0_bits_raddress : _GEN_447; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_entryid = io_in_0_valid ? io_in_0_bits_entryid : _GEN_446; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_arid = io_in_0_valid ? io_in_0_bits_arid : _GEN_445; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_ardata = io_in_0_valid ? io_in_0_bits_ardata : _GEN_444; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_respStatus = io_in_0_valid ? io_in_0_bits_respStatus : _GEN_442; // @[Arbiter.scala 141:26 143:19]
  assign io_out_bits_rsize = io_in_0_valid ? io_in_0_bits_rsize : _GEN_441; // @[Arbiter.scala 141:26 143:19]
  assign io_chosen = io_in_0_valid ? 5'h0 : _GEN_435; // @[Arbiter.scala 141:26 142:17]
endmodule
module ReadStack(
  input          clock,
  input          reset,
  output         io_axiReq_in_ar_ready,
  input          io_axiReq_in_ar_valid,
  input  [13:0]  io_axiReq_in_ar_bits_id,
  input  [34:0]  io_axiReq_in_ar_bits_addr,
  input  [7:0]   io_axiReq_in_ar_bits_len,
  input  [2:0]   io_axiReq_in_ar_bits_size,
  input  [1:0]   io_axiReq_in_ar_bits_burst,
  input          io_axiReq_in_ar_bits_lock,
  input  [3:0]   io_axiReq_in_ar_bits_cache,
  input  [2:0]   io_axiReq_in_ar_bits_prot,
  input  [3:0]   io_axiReq_in_ar_bits_qos,
  output         io_tlResp_in_d_ready,
  input          io_tlResp_in_d_valid,
  input  [2:0]   io_tlResp_in_d_bits_opcode,
  input  [1:0]   io_tlResp_in_d_bits_param,
  input  [2:0]   io_tlResp_in_d_bits_size,
  input  [18:0]  io_tlResp_in_d_bits_source,
  input  [4:0]   io_tlResp_in_d_bits_sink,
  input          io_tlResp_in_d_bits_denied,
  input  [255:0] io_tlResp_in_d_bits_data,
  input          io_tlResp_in_d_bits_corrupt,
  input          io_tlReq_out_a_ready,
  output         io_tlReq_out_a_valid,
  output [2:0]   io_tlReq_out_a_bits_opcode,
  output [2:0]   io_tlReq_out_a_bits_param,
  output [2:0]   io_tlReq_out_a_bits_size,
  output [18:0]  io_tlReq_out_a_bits_source,
  output [34:0]  io_tlReq_out_a_bits_address,
  output [31:0]  io_tlReq_out_a_bits_mask,
  output [255:0] io_tlReq_out_a_bits_data,
  output         io_tlReq_out_a_bits_corrupt,
  input          io_axiResp_out_r_ready,
  output         io_axiResp_out_r_valid,
  output [13:0]  io_axiResp_out_r_bits_id,
  output [255:0] io_axiResp_out_r_bits_data,
  output [1:0]   io_axiResp_out_r_bits_resp,
  output         io_axiResp_out_r_bits_last
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [255:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [255:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [255:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [255:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [63:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [255:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [63:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [255:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [63:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [255:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [63:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [255:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [63:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [255:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [63:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [255:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [63:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [255:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [63:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [255:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [63:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [255:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [63:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [255:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [63:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [255:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [63:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [255:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [63:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [255:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [63:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [255:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [63:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [255:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [63:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [255:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [63:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
  reg [255:0] _RAND_204;
  reg [31:0] _RAND_205;
  reg [31:0] _RAND_206;
  reg [31:0] _RAND_207;
  reg [31:0] _RAND_208;
  reg [31:0] _RAND_209;
  reg [31:0] _RAND_210;
  reg [63:0] _RAND_211;
  reg [31:0] _RAND_212;
  reg [31:0] _RAND_213;
  reg [255:0] _RAND_214;
  reg [31:0] _RAND_215;
  reg [31:0] _RAND_216;
  reg [31:0] _RAND_217;
  reg [31:0] _RAND_218;
  reg [31:0] _RAND_219;
  reg [31:0] _RAND_220;
  reg [63:0] _RAND_221;
  reg [31:0] _RAND_222;
  reg [31:0] _RAND_223;
  reg [255:0] _RAND_224;
  reg [31:0] _RAND_225;
  reg [31:0] _RAND_226;
  reg [31:0] _RAND_227;
  reg [31:0] _RAND_228;
  reg [31:0] _RAND_229;
  reg [31:0] _RAND_230;
  reg [63:0] _RAND_231;
  reg [31:0] _RAND_232;
  reg [31:0] _RAND_233;
  reg [255:0] _RAND_234;
  reg [31:0] _RAND_235;
  reg [31:0] _RAND_236;
  reg [31:0] _RAND_237;
  reg [31:0] _RAND_238;
  reg [31:0] _RAND_239;
  reg [31:0] _RAND_240;
  reg [63:0] _RAND_241;
  reg [31:0] _RAND_242;
  reg [31:0] _RAND_243;
  reg [255:0] _RAND_244;
  reg [31:0] _RAND_245;
  reg [31:0] _RAND_246;
  reg [31:0] _RAND_247;
  reg [31:0] _RAND_248;
  reg [31:0] _RAND_249;
  reg [31:0] _RAND_250;
  reg [63:0] _RAND_251;
  reg [31:0] _RAND_252;
  reg [31:0] _RAND_253;
  reg [255:0] _RAND_254;
  reg [31:0] _RAND_255;
  reg [31:0] _RAND_256;
  reg [31:0] _RAND_257;
  reg [31:0] _RAND_258;
  reg [31:0] _RAND_259;
  reg [31:0] _RAND_260;
  reg [63:0] _RAND_261;
  reg [31:0] _RAND_262;
  reg [31:0] _RAND_263;
  reg [255:0] _RAND_264;
  reg [31:0] _RAND_265;
  reg [31:0] _RAND_266;
  reg [31:0] _RAND_267;
  reg [31:0] _RAND_268;
  reg [31:0] _RAND_269;
  reg [31:0] _RAND_270;
  reg [63:0] _RAND_271;
  reg [31:0] _RAND_272;
  reg [31:0] _RAND_273;
  reg [255:0] _RAND_274;
  reg [31:0] _RAND_275;
  reg [31:0] _RAND_276;
  reg [31:0] _RAND_277;
  reg [31:0] _RAND_278;
  reg [31:0] _RAND_279;
  reg [31:0] _RAND_280;
  reg [63:0] _RAND_281;
  reg [31:0] _RAND_282;
  reg [31:0] _RAND_283;
  reg [255:0] _RAND_284;
  reg [31:0] _RAND_285;
  reg [31:0] _RAND_286;
  reg [31:0] _RAND_287;
  reg [31:0] _RAND_288;
  reg [31:0] _RAND_289;
  reg [31:0] _RAND_290;
  reg [63:0] _RAND_291;
  reg [31:0] _RAND_292;
  reg [31:0] _RAND_293;
  reg [255:0] _RAND_294;
  reg [31:0] _RAND_295;
  reg [31:0] _RAND_296;
  reg [31:0] _RAND_297;
  reg [31:0] _RAND_298;
  reg [31:0] _RAND_299;
  reg [31:0] _RAND_300;
  reg [63:0] _RAND_301;
  reg [31:0] _RAND_302;
  reg [31:0] _RAND_303;
  reg [255:0] _RAND_304;
  reg [31:0] _RAND_305;
  reg [31:0] _RAND_306;
  reg [31:0] _RAND_307;
  reg [31:0] _RAND_308;
  reg [31:0] _RAND_309;
  reg [31:0] _RAND_310;
  reg [63:0] _RAND_311;
  reg [31:0] _RAND_312;
  reg [31:0] _RAND_313;
  reg [255:0] _RAND_314;
  reg [31:0] _RAND_315;
  reg [31:0] _RAND_316;
  reg [31:0] _RAND_317;
  reg [31:0] _RAND_318;
  reg [31:0] _RAND_319;
`endif // RANDOMIZE_REG_INIT
  wire  axireqArb_io_in_0_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_0_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_0_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_0_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_0_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_0_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_0_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_1_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_1_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_1_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_1_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_1_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_1_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_1_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_2_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_2_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_2_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_2_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_2_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_2_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_2_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_3_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_3_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_3_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_3_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_3_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_3_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_3_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_4_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_4_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_4_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_4_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_4_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_4_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_4_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_5_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_5_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_5_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_5_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_5_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_5_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_5_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_6_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_6_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_6_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_6_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_6_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_6_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_6_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_7_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_7_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_7_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_7_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_7_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_7_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_7_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_8_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_8_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_8_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_8_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_8_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_8_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_8_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_9_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_9_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_9_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_9_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_9_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_9_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_9_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_10_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_10_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_10_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_10_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_10_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_10_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_10_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_11_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_11_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_11_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_11_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_11_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_11_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_11_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_12_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_12_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_12_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_12_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_12_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_12_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_12_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_13_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_13_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_13_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_13_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_13_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_13_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_13_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_14_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_14_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_14_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_14_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_14_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_14_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_14_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_15_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_15_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_15_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_15_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_15_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_15_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_15_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_16_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_16_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_16_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_16_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_16_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_16_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_16_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_17_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_17_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_17_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_17_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_17_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_17_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_17_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_18_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_18_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_18_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_18_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_18_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_18_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_18_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_19_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_19_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_19_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_19_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_19_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_19_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_19_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_20_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_20_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_20_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_20_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_20_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_20_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_20_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_21_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_21_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_21_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_21_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_21_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_21_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_21_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_22_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_22_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_22_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_22_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_22_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_22_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_22_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_23_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_23_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_23_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_23_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_23_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_23_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_23_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_24_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_24_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_24_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_24_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_24_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_24_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_24_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_25_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_25_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_25_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_25_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_25_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_25_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_25_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_26_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_26_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_26_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_26_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_26_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_26_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_26_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_27_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_27_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_27_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_27_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_27_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_27_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_27_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_28_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_28_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_28_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_28_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_28_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_28_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_28_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_29_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_29_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_29_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_29_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_29_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_29_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_29_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_30_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_30_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_30_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_30_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_30_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_30_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_30_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_in_31_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_in_31_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_in_31_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_in_31_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_in_31_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_in_31_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_in_31_bits_rsize; // @[ReadStack.scala 65:25]
  wire  axireqArb_io_out_valid; // @[ReadStack.scala 65:25]
  wire [34:0] axireqArb_io_out_bits_raddress; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_out_bits_entryid; // @[ReadStack.scala 65:25]
  wire [13:0] axireqArb_io_out_bits_arid; // @[ReadStack.scala 65:25]
  wire [255:0] axireqArb_io_out_bits_ardata; // @[ReadStack.scala 65:25]
  wire [3:0] axireqArb_io_out_bits_respStatus; // @[ReadStack.scala 65:25]
  wire [7:0] axireqArb_io_out_bits_rsize; // @[ReadStack.scala 65:25]
  wire [4:0] axireqArb_io_chosen; // @[ReadStack.scala 65:25]
  wire  axirespArb_io_in_0_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_0_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_0_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_0_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_0_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_0_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_0_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_1_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_1_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_1_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_1_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_1_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_1_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_1_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_2_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_2_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_2_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_2_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_2_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_2_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_2_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_3_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_3_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_3_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_3_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_3_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_3_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_3_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_4_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_4_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_4_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_4_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_4_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_4_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_4_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_5_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_5_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_5_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_5_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_5_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_5_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_5_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_6_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_6_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_6_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_6_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_6_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_6_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_6_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_7_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_7_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_7_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_7_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_7_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_7_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_7_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_8_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_8_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_8_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_8_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_8_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_8_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_8_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_9_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_9_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_9_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_9_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_9_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_9_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_9_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_10_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_10_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_10_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_10_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_10_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_10_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_10_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_11_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_11_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_11_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_11_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_11_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_11_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_11_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_12_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_12_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_12_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_12_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_12_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_12_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_12_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_13_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_13_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_13_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_13_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_13_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_13_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_13_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_14_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_14_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_14_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_14_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_14_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_14_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_14_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_15_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_15_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_15_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_15_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_15_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_15_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_15_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_16_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_16_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_16_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_16_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_16_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_16_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_16_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_17_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_17_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_17_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_17_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_17_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_17_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_17_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_18_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_18_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_18_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_18_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_18_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_18_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_18_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_19_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_19_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_19_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_19_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_19_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_19_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_19_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_20_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_20_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_20_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_20_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_20_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_20_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_20_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_21_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_21_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_21_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_21_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_21_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_21_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_21_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_22_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_22_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_22_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_22_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_22_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_22_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_22_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_23_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_23_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_23_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_23_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_23_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_23_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_23_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_24_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_24_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_24_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_24_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_24_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_24_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_24_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_25_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_25_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_25_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_25_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_25_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_25_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_25_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_26_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_26_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_26_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_26_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_26_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_26_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_26_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_27_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_27_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_27_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_27_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_27_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_27_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_27_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_28_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_28_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_28_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_28_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_28_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_28_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_28_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_29_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_29_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_29_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_29_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_29_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_29_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_29_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_30_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_30_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_30_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_30_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_30_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_30_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_30_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_in_31_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_in_31_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_in_31_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_in_31_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_in_31_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_in_31_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_in_31_bits_rsize; // @[ReadStack.scala 66:26]
  wire  axirespArb_io_out_valid; // @[ReadStack.scala 66:26]
  wire [34:0] axirespArb_io_out_bits_raddress; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_out_bits_entryid; // @[ReadStack.scala 66:26]
  wire [13:0] axirespArb_io_out_bits_arid; // @[ReadStack.scala 66:26]
  wire [255:0] axirespArb_io_out_bits_ardata; // @[ReadStack.scala 66:26]
  wire [3:0] axirespArb_io_out_bits_respStatus; // @[ReadStack.scala 66:26]
  wire [7:0] axirespArb_io_out_bits_rsize; // @[ReadStack.scala 66:26]
  wire [4:0] axirespArb_io_chosen; // @[ReadStack.scala 66:26]
  reg  readStack_0_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_0_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_0_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_0_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_0_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_0_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_0_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_0_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_0_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_0_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_1_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_1_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_1_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_1_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_1_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_1_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_1_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_1_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_1_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_1_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_2_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_2_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_2_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_2_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_2_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_2_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_2_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_2_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_2_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_2_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_3_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_3_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_3_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_3_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_3_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_3_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_3_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_3_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_3_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_3_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_4_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_4_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_4_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_4_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_4_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_4_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_4_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_4_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_4_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_4_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_5_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_5_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_5_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_5_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_5_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_5_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_5_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_5_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_5_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_5_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_6_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_6_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_6_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_6_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_6_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_6_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_6_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_6_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_6_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_6_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_7_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_7_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_7_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_7_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_7_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_7_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_7_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_7_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_7_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_7_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_8_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_8_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_8_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_8_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_8_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_8_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_8_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_8_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_8_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_8_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_9_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_9_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_9_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_9_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_9_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_9_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_9_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_9_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_9_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_9_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_10_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_10_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_10_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_10_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_10_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_10_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_10_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_10_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_10_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_10_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_11_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_11_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_11_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_11_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_11_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_11_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_11_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_11_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_11_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_11_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_12_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_12_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_12_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_12_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_12_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_12_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_12_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_12_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_12_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_12_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_13_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_13_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_13_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_13_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_13_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_13_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_13_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_13_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_13_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_13_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_14_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_14_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_14_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_14_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_14_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_14_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_14_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_14_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_14_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_14_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_15_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_15_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_15_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_15_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_15_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_15_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_15_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_15_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_15_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_15_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_16_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_16_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_16_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_16_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_16_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_16_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_16_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_16_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_16_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_16_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_17_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_17_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_17_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_17_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_17_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_17_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_17_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_17_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_17_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_17_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_18_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_18_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_18_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_18_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_18_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_18_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_18_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_18_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_18_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_18_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_19_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_19_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_19_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_19_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_19_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_19_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_19_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_19_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_19_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_19_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_20_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_20_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_20_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_20_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_20_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_20_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_20_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_20_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_20_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_20_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_21_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_21_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_21_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_21_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_21_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_21_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_21_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_21_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_21_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_21_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_22_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_22_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_22_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_22_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_22_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_22_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_22_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_22_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_22_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_22_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_23_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_23_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_23_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_23_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_23_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_23_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_23_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_23_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_23_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_23_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_24_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_24_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_24_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_24_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_24_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_24_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_24_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_24_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_24_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_24_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_25_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_25_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_25_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_25_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_25_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_25_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_25_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_25_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_25_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_25_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_26_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_26_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_26_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_26_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_26_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_26_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_26_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_26_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_26_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_26_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_27_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_27_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_27_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_27_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_27_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_27_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_27_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_27_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_27_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_27_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_28_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_28_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_28_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_28_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_28_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_28_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_28_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_28_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_28_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_28_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_29_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_29_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_29_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_29_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_29_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_29_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_29_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_29_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_29_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_29_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_30_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_30_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_30_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_30_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_30_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_30_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_30_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_30_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_30_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_30_BeatFifoId; // @[ReadStack.scala 63:26]
  reg  readStack_31_rvalid; // @[ReadStack.scala 63:26]
  reg [34:0] readStack_31_raddress; // @[ReadStack.scala 63:26]
  reg [4:0] readStack_31_entryid; // @[ReadStack.scala 63:26]
  reg [13:0] readStack_31_arid; // @[ReadStack.scala 63:26]
  reg [255:0] readStack_31_ardata; // @[ReadStack.scala 63:26]
  reg [1:0] readStack_31_readStatus; // @[ReadStack.scala 63:26]
  reg [3:0] readStack_31_respStatus; // @[ReadStack.scala 63:26]
  reg [7:0] readStack_31_rsize; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_31_entryFifoId; // @[ReadStack.scala 63:26]
  reg [5:0] readStack_31_BeatFifoId; // @[ReadStack.scala 63:26]
  wire [7:0] full_lo_lo = {readStack_24_rvalid,readStack_25_rvalid,readStack_26_rvalid,readStack_27_rvalid,
    readStack_28_rvalid,readStack_29_rvalid,readStack_30_rvalid,readStack_31_rvalid}; // @[Cat.scala 31:58]
  wire [15:0] full_lo = {readStack_16_rvalid,readStack_17_rvalid,readStack_18_rvalid,readStack_19_rvalid,
    readStack_20_rvalid,readStack_21_rvalid,readStack_22_rvalid,readStack_23_rvalid,full_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] full_hi_lo = {readStack_8_rvalid,readStack_9_rvalid,readStack_10_rvalid,readStack_11_rvalid,
    readStack_12_rvalid,readStack_13_rvalid,readStack_14_rvalid,readStack_15_rvalid}; // @[Cat.scala 31:58]
  wire [31:0] _full_T = {readStack_0_rvalid,readStack_1_rvalid,readStack_2_rvalid,readStack_3_rvalid,readStack_4_rvalid,
    readStack_5_rvalid,readStack_6_rvalid,readStack_7_rvalid,full_hi_lo,full_lo}; // @[Cat.scala 31:58]
  wire  full = &_full_T; // @[ReadStack.scala 69:43]
  wire  alloc = ~full & io_axiReq_in_ar_valid; // @[ReadStack.scala 70:21]
  wire  _idxInsert_T = ~readStack_0_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_1 = ~readStack_1_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_2 = ~readStack_2_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_3 = ~readStack_3_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_4 = ~readStack_4_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_5 = ~readStack_5_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_6 = ~readStack_6_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_7 = ~readStack_7_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_8 = ~readStack_8_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_9 = ~readStack_9_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_10 = ~readStack_10_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_11 = ~readStack_11_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_12 = ~readStack_12_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_13 = ~readStack_13_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_14 = ~readStack_14_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_15 = ~readStack_15_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_16 = ~readStack_16_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_17 = ~readStack_17_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_18 = ~readStack_18_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_19 = ~readStack_19_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_20 = ~readStack_20_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_21 = ~readStack_21_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_22 = ~readStack_22_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_23 = ~readStack_23_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_24 = ~readStack_24_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_25 = ~readStack_25_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_26 = ~readStack_26_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_27 = ~readStack_27_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_28 = ~readStack_28_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_29 = ~readStack_29_rvalid; // @[ReadStack.scala 74:59]
  wire  _idxInsert_T_30 = ~readStack_30_rvalid; // @[ReadStack.scala 74:59]
  wire [4:0] _idxInsert_T_32 = _idxInsert_T_30 ? 5'h1e : 5'h1f; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_33 = _idxInsert_T_29 ? 5'h1d : _idxInsert_T_32; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_34 = _idxInsert_T_28 ? 5'h1c : _idxInsert_T_33; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_35 = _idxInsert_T_27 ? 5'h1b : _idxInsert_T_34; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_36 = _idxInsert_T_26 ? 5'h1a : _idxInsert_T_35; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_37 = _idxInsert_T_25 ? 5'h19 : _idxInsert_T_36; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_38 = _idxInsert_T_24 ? 5'h18 : _idxInsert_T_37; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_39 = _idxInsert_T_23 ? 5'h17 : _idxInsert_T_38; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_40 = _idxInsert_T_22 ? 5'h16 : _idxInsert_T_39; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_41 = _idxInsert_T_21 ? 5'h15 : _idxInsert_T_40; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_42 = _idxInsert_T_20 ? 5'h14 : _idxInsert_T_41; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_43 = _idxInsert_T_19 ? 5'h13 : _idxInsert_T_42; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_44 = _idxInsert_T_18 ? 5'h12 : _idxInsert_T_43; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_45 = _idxInsert_T_17 ? 5'h11 : _idxInsert_T_44; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_46 = _idxInsert_T_16 ? 5'h10 : _idxInsert_T_45; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_47 = _idxInsert_T_15 ? 5'hf : _idxInsert_T_46; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_48 = _idxInsert_T_14 ? 5'he : _idxInsert_T_47; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_49 = _idxInsert_T_13 ? 5'hd : _idxInsert_T_48; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_50 = _idxInsert_T_12 ? 5'hc : _idxInsert_T_49; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_51 = _idxInsert_T_11 ? 5'hb : _idxInsert_T_50; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_52 = _idxInsert_T_10 ? 5'ha : _idxInsert_T_51; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_53 = _idxInsert_T_9 ? 5'h9 : _idxInsert_T_52; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_54 = _idxInsert_T_8 ? 5'h8 : _idxInsert_T_53; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_55 = _idxInsert_T_7 ? 5'h7 : _idxInsert_T_54; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_56 = _idxInsert_T_6 ? 5'h6 : _idxInsert_T_55; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_57 = _idxInsert_T_5 ? 5'h5 : _idxInsert_T_56; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_58 = _idxInsert_T_4 ? 5'h4 : _idxInsert_T_57; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_59 = _idxInsert_T_3 ? 5'h3 : _idxInsert_T_58; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_60 = _idxInsert_T_2 ? 5'h2 : _idxInsert_T_59; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_61 = _idxInsert_T_1 ? 5'h1 : _idxInsert_T_60; // @[Mux.scala 47:70]
  wire [4:0] _idxInsert_T_62 = _idxInsert_T ? 5'h0 : _idxInsert_T_61; // @[Mux.scala 47:70]
  wire [4:0] idxInsert = alloc ? _idxInsert_T_62 : 5'h0; // @[ReadStack.scala 74:22]
  wire [15:0] _r_size1_T = {io_axiReq_in_ar_bits_len,8'hff}; // @[Cat.scala 31:58]
  wire [22:0] _GEN_544 = {{7'd0}, _r_size1_T}; // @[Bundles.scala 34:21]
  wire [22:0] _r_size1_T_1 = _GEN_544 << io_axiReq_in_ar_bits_size; // @[Bundles.scala 34:21]
  wire [14:0] r_size1 = _r_size1_T_1[22:8]; // @[Bundles.scala 34:30]
  wire  _GEN_0 = 5'h0 == idxInsert | readStack_0_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_1 = 5'h1 == idxInsert | readStack_1_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_2 = 5'h2 == idxInsert | readStack_2_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_3 = 5'h3 == idxInsert | readStack_3_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_4 = 5'h4 == idxInsert | readStack_4_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_5 = 5'h5 == idxInsert | readStack_5_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_6 = 5'h6 == idxInsert | readStack_6_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_7 = 5'h7 == idxInsert | readStack_7_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_8 = 5'h8 == idxInsert | readStack_8_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_9 = 5'h9 == idxInsert | readStack_9_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_10 = 5'ha == idxInsert | readStack_10_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_11 = 5'hb == idxInsert | readStack_11_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_12 = 5'hc == idxInsert | readStack_12_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_13 = 5'hd == idxInsert | readStack_13_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_14 = 5'he == idxInsert | readStack_14_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_15 = 5'hf == idxInsert | readStack_15_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_16 = 5'h10 == idxInsert | readStack_16_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_17 = 5'h11 == idxInsert | readStack_17_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_18 = 5'h12 == idxInsert | readStack_18_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_19 = 5'h13 == idxInsert | readStack_19_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_20 = 5'h14 == idxInsert | readStack_20_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_21 = 5'h15 == idxInsert | readStack_21_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_22 = 5'h16 == idxInsert | readStack_22_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_23 = 5'h17 == idxInsert | readStack_23_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_24 = 5'h18 == idxInsert | readStack_24_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_25 = 5'h19 == idxInsert | readStack_25_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_26 = 5'h1a == idxInsert | readStack_26_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_27 = 5'h1b == idxInsert | readStack_27_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_28 = 5'h1c == idxInsert | readStack_28_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_29 = 5'h1d == idxInsert | readStack_29_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_30 = 5'h1e == idxInsert | readStack_30_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire  _GEN_31 = 5'h1f == idxInsert | readStack_31_rvalid; // @[ReadStack.scala 83:{20,20} 63:26]
  wire [1:0] _GEN_128 = 5'h0 == idxInsert ? 2'h1 : readStack_0_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_129 = 5'h1 == idxInsert ? 2'h1 : readStack_1_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_130 = 5'h2 == idxInsert ? 2'h1 : readStack_2_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_131 = 5'h3 == idxInsert ? 2'h1 : readStack_3_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_132 = 5'h4 == idxInsert ? 2'h1 : readStack_4_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_133 = 5'h5 == idxInsert ? 2'h1 : readStack_5_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_134 = 5'h6 == idxInsert ? 2'h1 : readStack_6_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_135 = 5'h7 == idxInsert ? 2'h1 : readStack_7_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_136 = 5'h8 == idxInsert ? 2'h1 : readStack_8_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_137 = 5'h9 == idxInsert ? 2'h1 : readStack_9_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_138 = 5'ha == idxInsert ? 2'h1 : readStack_10_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_139 = 5'hb == idxInsert ? 2'h1 : readStack_11_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_140 = 5'hc == idxInsert ? 2'h1 : readStack_12_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_141 = 5'hd == idxInsert ? 2'h1 : readStack_13_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_142 = 5'he == idxInsert ? 2'h1 : readStack_14_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_143 = 5'hf == idxInsert ? 2'h1 : readStack_15_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_144 = 5'h10 == idxInsert ? 2'h1 : readStack_16_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_145 = 5'h11 == idxInsert ? 2'h1 : readStack_17_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_146 = 5'h12 == idxInsert ? 2'h1 : readStack_18_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_147 = 5'h13 == idxInsert ? 2'h1 : readStack_19_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_148 = 5'h14 == idxInsert ? 2'h1 : readStack_20_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_149 = 5'h15 == idxInsert ? 2'h1 : readStack_21_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_150 = 5'h16 == idxInsert ? 2'h1 : readStack_22_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_151 = 5'h17 == idxInsert ? 2'h1 : readStack_23_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_152 = 5'h18 == idxInsert ? 2'h1 : readStack_24_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_153 = 5'h19 == idxInsert ? 2'h1 : readStack_25_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_154 = 5'h1a == idxInsert ? 2'h1 : readStack_26_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_155 = 5'h1b == idxInsert ? 2'h1 : readStack_27_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_156 = 5'h1c == idxInsert ? 2'h1 : readStack_28_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_157 = 5'h1d == idxInsert ? 2'h1 : readStack_29_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_158 = 5'h1e == idxInsert ? 2'h1 : readStack_30_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire [1:0] _GEN_159 = 5'h1f == idxInsert ? 2'h1 : readStack_31_readStatus; // @[ReadStack.scala 87:{24,24} 63:26]
  wire  _GEN_192 = alloc ? _GEN_0 : readStack_0_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_193 = alloc ? _GEN_1 : readStack_1_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_194 = alloc ? _GEN_2 : readStack_2_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_195 = alloc ? _GEN_3 : readStack_3_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_196 = alloc ? _GEN_4 : readStack_4_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_197 = alloc ? _GEN_5 : readStack_5_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_198 = alloc ? _GEN_6 : readStack_6_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_199 = alloc ? _GEN_7 : readStack_7_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_200 = alloc ? _GEN_8 : readStack_8_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_201 = alloc ? _GEN_9 : readStack_9_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_202 = alloc ? _GEN_10 : readStack_10_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_203 = alloc ? _GEN_11 : readStack_11_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_204 = alloc ? _GEN_12 : readStack_12_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_205 = alloc ? _GEN_13 : readStack_13_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_206 = alloc ? _GEN_14 : readStack_14_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_207 = alloc ? _GEN_15 : readStack_15_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_208 = alloc ? _GEN_16 : readStack_16_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_209 = alloc ? _GEN_17 : readStack_17_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_210 = alloc ? _GEN_18 : readStack_18_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_211 = alloc ? _GEN_19 : readStack_19_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_212 = alloc ? _GEN_20 : readStack_20_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_213 = alloc ? _GEN_21 : readStack_21_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_214 = alloc ? _GEN_22 : readStack_22_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_215 = alloc ? _GEN_23 : readStack_23_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_216 = alloc ? _GEN_24 : readStack_24_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_217 = alloc ? _GEN_25 : readStack_25_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_218 = alloc ? _GEN_26 : readStack_26_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_219 = alloc ? _GEN_27 : readStack_27_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_220 = alloc ? _GEN_28 : readStack_28_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_221 = alloc ? _GEN_29 : readStack_29_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_222 = alloc ? _GEN_30 : readStack_30_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire  _GEN_223 = alloc ? _GEN_31 : readStack_31_rvalid; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_320 = alloc ? _GEN_128 : readStack_0_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_321 = alloc ? _GEN_129 : readStack_1_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_322 = alloc ? _GEN_130 : readStack_2_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_323 = alloc ? _GEN_131 : readStack_3_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_324 = alloc ? _GEN_132 : readStack_4_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_325 = alloc ? _GEN_133 : readStack_5_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_326 = alloc ? _GEN_134 : readStack_6_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_327 = alloc ? _GEN_135 : readStack_7_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_328 = alloc ? _GEN_136 : readStack_8_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_329 = alloc ? _GEN_137 : readStack_9_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_330 = alloc ? _GEN_138 : readStack_10_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_331 = alloc ? _GEN_139 : readStack_11_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_332 = alloc ? _GEN_140 : readStack_12_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_333 = alloc ? _GEN_141 : readStack_13_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_334 = alloc ? _GEN_142 : readStack_14_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_335 = alloc ? _GEN_143 : readStack_15_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_336 = alloc ? _GEN_144 : readStack_16_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_337 = alloc ? _GEN_145 : readStack_17_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_338 = alloc ? _GEN_146 : readStack_18_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_339 = alloc ? _GEN_147 : readStack_19_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_340 = alloc ? _GEN_148 : readStack_20_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_341 = alloc ? _GEN_149 : readStack_21_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_342 = alloc ? _GEN_150 : readStack_22_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_343 = alloc ? _GEN_151 : readStack_23_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_344 = alloc ? _GEN_152 : readStack_24_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_345 = alloc ? _GEN_153 : readStack_25_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_346 = alloc ? _GEN_154 : readStack_26_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_347 = alloc ? _GEN_155 : readStack_27_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_348 = alloc ? _GEN_156 : readStack_28_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_349 = alloc ? _GEN_157 : readStack_29_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_350 = alloc ? _GEN_158 : readStack_30_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [1:0] _GEN_351 = alloc ? _GEN_159 : readStack_31_readStatus; // @[ReadStack.scala 63:26 78:5]
  wire [2:0] _GEN_1184 = {{1'd0}, readStack_0_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T = _GEN_1184 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1185 = {{1'd0}, readStack_1_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_1 = _GEN_1185 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1186 = {{1'd0}, readStack_2_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_2 = _GEN_1186 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1187 = {{1'd0}, readStack_3_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_3 = _GEN_1187 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1188 = {{1'd0}, readStack_4_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_4 = _GEN_1188 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1189 = {{1'd0}, readStack_5_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_5 = _GEN_1189 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1190 = {{1'd0}, readStack_6_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_6 = _GEN_1190 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1191 = {{1'd0}, readStack_7_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_7 = _GEN_1191 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1192 = {{1'd0}, readStack_8_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_8 = _GEN_1192 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1193 = {{1'd0}, readStack_9_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_9 = _GEN_1193 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1194 = {{1'd0}, readStack_10_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_10 = _GEN_1194 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1195 = {{1'd0}, readStack_11_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_11 = _GEN_1195 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1196 = {{1'd0}, readStack_12_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_12 = _GEN_1196 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1197 = {{1'd0}, readStack_13_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_13 = _GEN_1197 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1198 = {{1'd0}, readStack_14_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_14 = _GEN_1198 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1199 = {{1'd0}, readStack_15_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_15 = _GEN_1199 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1200 = {{1'd0}, readStack_16_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_16 = _GEN_1200 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1201 = {{1'd0}, readStack_17_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_17 = _GEN_1201 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1202 = {{1'd0}, readStack_18_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_18 = _GEN_1202 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1203 = {{1'd0}, readStack_19_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_19 = _GEN_1203 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1204 = {{1'd0}, readStack_20_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_20 = _GEN_1204 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1205 = {{1'd0}, readStack_21_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_21 = _GEN_1205 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1206 = {{1'd0}, readStack_22_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_22 = _GEN_1206 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1207 = {{1'd0}, readStack_23_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_23 = _GEN_1207 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1208 = {{1'd0}, readStack_24_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_24 = _GEN_1208 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1209 = {{1'd0}, readStack_25_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_25 = _GEN_1209 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1210 = {{1'd0}, readStack_26_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_26 = _GEN_1210 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1211 = {{1'd0}, readStack_27_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_27 = _GEN_1211 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1212 = {{1'd0}, readStack_28_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_28 = _GEN_1212 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1213 = {{1'd0}, readStack_29_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_29 = _GEN_1213 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1214 = {{1'd0}, readStack_30_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_30 = _GEN_1214 == 3'h1; // @[ReadStack.scala 98:53]
  wire [2:0] _GEN_1215 = {{1'd0}, readStack_31_readStatus}; // @[ReadStack.scala 98:53]
  wire  _hasWaitTLReq_T_31 = _GEN_1215 == 3'h1; // @[ReadStack.scala 98:53]
  wire  _axireqArb_io_in_0_valid_T_1 = readStack_0_rvalid & _hasWaitTLReq_T; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_1_valid_T_1 = readStack_1_rvalid & _hasWaitTLReq_T_1; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_2_valid_T_1 = readStack_2_rvalid & _hasWaitTLReq_T_2; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_3_valid_T_1 = readStack_3_rvalid & _hasWaitTLReq_T_3; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_4_valid_T_1 = readStack_4_rvalid & _hasWaitTLReq_T_4; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_5_valid_T_1 = readStack_5_rvalid & _hasWaitTLReq_T_5; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_6_valid_T_1 = readStack_6_rvalid & _hasWaitTLReq_T_6; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_7_valid_T_1 = readStack_7_rvalid & _hasWaitTLReq_T_7; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_8_valid_T_1 = readStack_8_rvalid & _hasWaitTLReq_T_8; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_9_valid_T_1 = readStack_9_rvalid & _hasWaitTLReq_T_9; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_10_valid_T_1 = readStack_10_rvalid & _hasWaitTLReq_T_10; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_11_valid_T_1 = readStack_11_rvalid & _hasWaitTLReq_T_11; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_12_valid_T_1 = readStack_12_rvalid & _hasWaitTLReq_T_12; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_13_valid_T_1 = readStack_13_rvalid & _hasWaitTLReq_T_13; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_14_valid_T_1 = readStack_14_rvalid & _hasWaitTLReq_T_14; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_15_valid_T_1 = readStack_15_rvalid & _hasWaitTLReq_T_15; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_16_valid_T_1 = readStack_16_rvalid & _hasWaitTLReq_T_16; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_17_valid_T_1 = readStack_17_rvalid & _hasWaitTLReq_T_17; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_18_valid_T_1 = readStack_18_rvalid & _hasWaitTLReq_T_18; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_19_valid_T_1 = readStack_19_rvalid & _hasWaitTLReq_T_19; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_20_valid_T_1 = readStack_20_rvalid & _hasWaitTLReq_T_20; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_21_valid_T_1 = readStack_21_rvalid & _hasWaitTLReq_T_21; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_22_valid_T_1 = readStack_22_rvalid & _hasWaitTLReq_T_22; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_23_valid_T_1 = readStack_23_rvalid & _hasWaitTLReq_T_23; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_24_valid_T_1 = readStack_24_rvalid & _hasWaitTLReq_T_24; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_25_valid_T_1 = readStack_25_rvalid & _hasWaitTLReq_T_25; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_26_valid_T_1 = readStack_26_rvalid & _hasWaitTLReq_T_26; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_27_valid_T_1 = readStack_27_rvalid & _hasWaitTLReq_T_27; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_28_valid_T_1 = readStack_28_rvalid & _hasWaitTLReq_T_28; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_29_valid_T_1 = readStack_29_rvalid & _hasWaitTLReq_T_29; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_30_valid_T_1 = readStack_30_rvalid & _hasWaitTLReq_T_30; // @[ReadStack.scala 104:28]
  wire  _axireqArb_io_in_31_valid_T_1 = readStack_31_rvalid & _hasWaitTLReq_T_31; // @[ReadStack.scala 104:28]
  wire [7:0] _io_tlReq_out_a_bits_mask_sizeOH_T = axireqArb_io_out_bits_rsize; // @[Misc.scala 201:34]
  wire [1:0] io_tlReq_out_a_bits_mask_sizeOH_shiftAmount = _io_tlReq_out_a_bits_mask_sizeOH_T[1:0]; // @[OneHot.scala 63:49]
  wire [3:0] _io_tlReq_out_a_bits_mask_sizeOH_T_1 = 4'h1 << io_tlReq_out_a_bits_mask_sizeOH_shiftAmount; // @[OneHot.scala 64:12]
  wire [2:0] io_tlReq_out_a_bits_mask_sizeOH = _io_tlReq_out_a_bits_mask_sizeOH_T_1[2:0] | 3'h1; // @[Misc.scala 201:81]
  wire  _io_tlReq_out_a_bits_mask_T = axireqArb_io_out_bits_rsize >= 8'h3; // @[Misc.scala 205:21]
  wire  io_tlReq_out_a_bits_mask_size = io_tlReq_out_a_bits_mask_sizeOH[2]; // @[Misc.scala 208:26]
  wire  io_tlReq_out_a_bits_mask_bit = axireqArb_io_out_bits_raddress[2]; // @[Misc.scala 209:26]
  wire  io_tlReq_out_a_bits_mask_nbit = ~io_tlReq_out_a_bits_mask_bit; // @[Misc.scala 210:20]
  wire  io_tlReq_out_a_bits_mask_acc = _io_tlReq_out_a_bits_mask_T | io_tlReq_out_a_bits_mask_size &
    io_tlReq_out_a_bits_mask_nbit; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_acc_1 = _io_tlReq_out_a_bits_mask_T | io_tlReq_out_a_bits_mask_size &
    io_tlReq_out_a_bits_mask_bit; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_size_1 = io_tlReq_out_a_bits_mask_sizeOH[1]; // @[Misc.scala 208:26]
  wire  io_tlReq_out_a_bits_mask_bit_1 = axireqArb_io_out_bits_raddress[1]; // @[Misc.scala 209:26]
  wire  io_tlReq_out_a_bits_mask_nbit_1 = ~io_tlReq_out_a_bits_mask_bit_1; // @[Misc.scala 210:20]
  wire  io_tlReq_out_a_bits_mask_eq_2 = io_tlReq_out_a_bits_mask_nbit & io_tlReq_out_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_2 = io_tlReq_out_a_bits_mask_acc | io_tlReq_out_a_bits_mask_size_1 &
    io_tlReq_out_a_bits_mask_eq_2; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_3 = io_tlReq_out_a_bits_mask_nbit & io_tlReq_out_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_3 = io_tlReq_out_a_bits_mask_acc | io_tlReq_out_a_bits_mask_size_1 &
    io_tlReq_out_a_bits_mask_eq_3; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_4 = io_tlReq_out_a_bits_mask_bit & io_tlReq_out_a_bits_mask_nbit_1; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_4 = io_tlReq_out_a_bits_mask_acc_1 | io_tlReq_out_a_bits_mask_size_1 &
    io_tlReq_out_a_bits_mask_eq_4; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_5 = io_tlReq_out_a_bits_mask_bit & io_tlReq_out_a_bits_mask_bit_1; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_5 = io_tlReq_out_a_bits_mask_acc_1 | io_tlReq_out_a_bits_mask_size_1 &
    io_tlReq_out_a_bits_mask_eq_5; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_size_2 = io_tlReq_out_a_bits_mask_sizeOH[0]; // @[Misc.scala 208:26]
  wire  io_tlReq_out_a_bits_mask_bit_2 = axireqArb_io_out_bits_raddress[0]; // @[Misc.scala 209:26]
  wire  io_tlReq_out_a_bits_mask_nbit_2 = ~io_tlReq_out_a_bits_mask_bit_2; // @[Misc.scala 210:20]
  wire  io_tlReq_out_a_bits_mask_eq_6 = io_tlReq_out_a_bits_mask_eq_2 & io_tlReq_out_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_6 = io_tlReq_out_a_bits_mask_acc_2 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_6; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_7 = io_tlReq_out_a_bits_mask_eq_2 & io_tlReq_out_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_7 = io_tlReq_out_a_bits_mask_acc_2 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_7; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_8 = io_tlReq_out_a_bits_mask_eq_3 & io_tlReq_out_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_8 = io_tlReq_out_a_bits_mask_acc_3 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_8; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_9 = io_tlReq_out_a_bits_mask_eq_3 & io_tlReq_out_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_9 = io_tlReq_out_a_bits_mask_acc_3 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_9; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_10 = io_tlReq_out_a_bits_mask_eq_4 & io_tlReq_out_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_10 = io_tlReq_out_a_bits_mask_acc_4 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_10; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_11 = io_tlReq_out_a_bits_mask_eq_4 & io_tlReq_out_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_11 = io_tlReq_out_a_bits_mask_acc_4 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_11; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_12 = io_tlReq_out_a_bits_mask_eq_5 & io_tlReq_out_a_bits_mask_nbit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_12 = io_tlReq_out_a_bits_mask_acc_5 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_12; // @[Misc.scala 214:29]
  wire  io_tlReq_out_a_bits_mask_eq_13 = io_tlReq_out_a_bits_mask_eq_5 & io_tlReq_out_a_bits_mask_bit_2; // @[Misc.scala 213:27]
  wire  io_tlReq_out_a_bits_mask_acc_13 = io_tlReq_out_a_bits_mask_acc_5 | io_tlReq_out_a_bits_mask_size_2 &
    io_tlReq_out_a_bits_mask_eq_13; // @[Misc.scala 214:29]
  wire [7:0] _io_tlReq_out_a_bits_mask_T_1 = {io_tlReq_out_a_bits_mask_acc_13,io_tlReq_out_a_bits_mask_acc_12,
    io_tlReq_out_a_bits_mask_acc_11,io_tlReq_out_a_bits_mask_acc_10,io_tlReq_out_a_bits_mask_acc_9,
    io_tlReq_out_a_bits_mask_acc_8,io_tlReq_out_a_bits_mask_acc_7,io_tlReq_out_a_bits_mask_acc_6}; // @[Cat.scala 31:58]
  wire  _T = io_axiReq_in_ar_ready & io_axiReq_in_ar_valid; // @[Decoupled.scala 50:35]
  wire  _T_1 = io_tlReq_out_a_ready & io_tlReq_out_a_valid; // @[Decoupled.scala 50:35]
  wire  _T_2 = _T & _T_1; // @[ReadStack.scala 126:29]
  wire [7:0] readStack_entryFifoId_lo_lo = {_axireqArb_io_in_24_valid_T_1,_axireqArb_io_in_25_valid_T_1,
    _axireqArb_io_in_26_valid_T_1,_axireqArb_io_in_27_valid_T_1,_axireqArb_io_in_28_valid_T_1,
    _axireqArb_io_in_29_valid_T_1,_axireqArb_io_in_30_valid_T_1,_axireqArb_io_in_31_valid_T_1}; // @[Cat.scala 31:58]
  wire [15:0] readStack_entryFifoId_lo = {_axireqArb_io_in_16_valid_T_1,_axireqArb_io_in_17_valid_T_1,
    _axireqArb_io_in_18_valid_T_1,_axireqArb_io_in_19_valid_T_1,_axireqArb_io_in_20_valid_T_1,
    _axireqArb_io_in_21_valid_T_1,_axireqArb_io_in_22_valid_T_1,_axireqArb_io_in_23_valid_T_1,
    readStack_entryFifoId_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] readStack_entryFifoId_hi_lo = {_axireqArb_io_in_8_valid_T_1,_axireqArb_io_in_9_valid_T_1,
    _axireqArb_io_in_10_valid_T_1,_axireqArb_io_in_11_valid_T_1,_axireqArb_io_in_12_valid_T_1,
    _axireqArb_io_in_13_valid_T_1,_axireqArb_io_in_14_valid_T_1,_axireqArb_io_in_15_valid_T_1}; // @[Cat.scala 31:58]
  wire [31:0] _readStack_entryFifoId_T_64 = {_axireqArb_io_in_0_valid_T_1,_axireqArb_io_in_1_valid_T_1,
    _axireqArb_io_in_2_valid_T_1,_axireqArb_io_in_3_valid_T_1,_axireqArb_io_in_4_valid_T_1,_axireqArb_io_in_5_valid_T_1,
    _axireqArb_io_in_6_valid_T_1,_axireqArb_io_in_7_valid_T_1,readStack_entryFifoId_hi_lo,readStack_entryFifoId_lo}; // @[Cat.scala 31:58]
  wire [1:0] _readStack_entryFifoId_T_97 = _readStack_entryFifoId_T_64[0] + _readStack_entryFifoId_T_64[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_99 = _readStack_entryFifoId_T_64[2] + _readStack_entryFifoId_T_64[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_101 = _readStack_entryFifoId_T_97 + _readStack_entryFifoId_T_99; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_103 = _readStack_entryFifoId_T_64[4] + _readStack_entryFifoId_T_64[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_105 = _readStack_entryFifoId_T_64[6] + _readStack_entryFifoId_T_64[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_107 = _readStack_entryFifoId_T_103 + _readStack_entryFifoId_T_105; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_entryFifoId_T_109 = _readStack_entryFifoId_T_101 + _readStack_entryFifoId_T_107; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_111 = _readStack_entryFifoId_T_64[8] + _readStack_entryFifoId_T_64[9]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_113 = _readStack_entryFifoId_T_64[10] + _readStack_entryFifoId_T_64[11]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_115 = _readStack_entryFifoId_T_111 + _readStack_entryFifoId_T_113; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_117 = _readStack_entryFifoId_T_64[12] + _readStack_entryFifoId_T_64[13]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_119 = _readStack_entryFifoId_T_64[14] + _readStack_entryFifoId_T_64[15]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_121 = _readStack_entryFifoId_T_117 + _readStack_entryFifoId_T_119; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_entryFifoId_T_123 = _readStack_entryFifoId_T_115 + _readStack_entryFifoId_T_121; // @[Bitwise.scala 48:55]
  wire [4:0] _readStack_entryFifoId_T_125 = _readStack_entryFifoId_T_109 + _readStack_entryFifoId_T_123; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_127 = _readStack_entryFifoId_T_64[16] + _readStack_entryFifoId_T_64[17]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_129 = _readStack_entryFifoId_T_64[18] + _readStack_entryFifoId_T_64[19]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_131 = _readStack_entryFifoId_T_127 + _readStack_entryFifoId_T_129; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_133 = _readStack_entryFifoId_T_64[20] + _readStack_entryFifoId_T_64[21]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_135 = _readStack_entryFifoId_T_64[22] + _readStack_entryFifoId_T_64[23]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_137 = _readStack_entryFifoId_T_133 + _readStack_entryFifoId_T_135; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_entryFifoId_T_139 = _readStack_entryFifoId_T_131 + _readStack_entryFifoId_T_137; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_141 = _readStack_entryFifoId_T_64[24] + _readStack_entryFifoId_T_64[25]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_143 = _readStack_entryFifoId_T_64[26] + _readStack_entryFifoId_T_64[27]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_145 = _readStack_entryFifoId_T_141 + _readStack_entryFifoId_T_143; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_147 = _readStack_entryFifoId_T_64[28] + _readStack_entryFifoId_T_64[29]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_entryFifoId_T_149 = _readStack_entryFifoId_T_64[30] + _readStack_entryFifoId_T_64[31]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_entryFifoId_T_151 = _readStack_entryFifoId_T_147 + _readStack_entryFifoId_T_149; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_entryFifoId_T_153 = _readStack_entryFifoId_T_145 + _readStack_entryFifoId_T_151; // @[Bitwise.scala 48:55]
  wire [4:0] _readStack_entryFifoId_T_155 = _readStack_entryFifoId_T_139 + _readStack_entryFifoId_T_153; // @[Bitwise.scala 48:55]
  wire [5:0] _readStack_entryFifoId_T_157 = _readStack_entryFifoId_T_125 + _readStack_entryFifoId_T_155; // @[Bitwise.scala 48:55]
  wire [5:0] _readStack_entryFifoId_T_160 = _readStack_entryFifoId_T_157 - 6'h1; // @[ReadStack.scala 130:105]
  wire [5:0] _GEN_384 = 5'h0 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_0_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_385 = 5'h1 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_1_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_386 = 5'h2 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_2_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_387 = 5'h3 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_3_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_388 = 5'h4 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_4_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_389 = 5'h5 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_5_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_390 = 5'h6 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_6_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_391 = 5'h7 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_7_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_392 = 5'h8 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_8_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_393 = 5'h9 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_9_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_394 = 5'ha == idxInsert ? _readStack_entryFifoId_T_160 : readStack_10_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_395 = 5'hb == idxInsert ? _readStack_entryFifoId_T_160 : readStack_11_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_396 = 5'hc == idxInsert ? _readStack_entryFifoId_T_160 : readStack_12_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_397 = 5'hd == idxInsert ? _readStack_entryFifoId_T_160 : readStack_13_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_398 = 5'he == idxInsert ? _readStack_entryFifoId_T_160 : readStack_14_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_399 = 5'hf == idxInsert ? _readStack_entryFifoId_T_160 : readStack_15_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_400 = 5'h10 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_16_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_401 = 5'h11 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_17_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_402 = 5'h12 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_18_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_403 = 5'h13 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_19_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_404 = 5'h14 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_20_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_405 = 5'h15 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_21_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_406 = 5'h16 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_22_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_407 = 5'h17 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_23_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_408 = 5'h18 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_24_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_409 = 5'h19 == idxInsert ? _readStack_entryFifoId_T_160 : readStack_25_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_410 = 5'h1a == idxInsert ? _readStack_entryFifoId_T_160 : readStack_26_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_411 = 5'h1b == idxInsert ? _readStack_entryFifoId_T_160 : readStack_27_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_412 = 5'h1c == idxInsert ? _readStack_entryFifoId_T_160 : readStack_28_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_413 = 5'h1d == idxInsert ? _readStack_entryFifoId_T_160 : readStack_29_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_414 = 5'h1e == idxInsert ? _readStack_entryFifoId_T_160 : readStack_30_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire [5:0] _GEN_415 = 5'h1f == idxInsert ? _readStack_entryFifoId_T_160 : readStack_31_entryFifoId; // @[ReadStack.scala 130:{27,27} 63:26]
  wire  _T_6 = _T & ~_T_1; // @[ReadStack.scala 131:37]
  wire [1:0] _readStack_entryFifoId_T_225 = _axireqArb_io_in_0_valid_T_1 + _axireqArb_io_in_1_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_227 = _axireqArb_io_in_2_valid_T_1 + _axireqArb_io_in_3_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_229 = _readStack_entryFifoId_T_225 + _readStack_entryFifoId_T_227; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_231 = _axireqArb_io_in_4_valid_T_1 + _axireqArb_io_in_5_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_233 = _axireqArb_io_in_6_valid_T_1 + _axireqArb_io_in_7_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_235 = _readStack_entryFifoId_T_231 + _readStack_entryFifoId_T_233; // @[ReadStack.scala 135:45]
  wire [3:0] _readStack_entryFifoId_T_237 = _readStack_entryFifoId_T_229 + _readStack_entryFifoId_T_235; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_239 = _axireqArb_io_in_8_valid_T_1 + _axireqArb_io_in_9_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_241 = _axireqArb_io_in_10_valid_T_1 + _axireqArb_io_in_11_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_243 = _readStack_entryFifoId_T_239 + _readStack_entryFifoId_T_241; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_245 = _axireqArb_io_in_12_valid_T_1 + _axireqArb_io_in_13_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_247 = _axireqArb_io_in_14_valid_T_1 + _axireqArb_io_in_15_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_249 = _readStack_entryFifoId_T_245 + _readStack_entryFifoId_T_247; // @[ReadStack.scala 135:45]
  wire [3:0] _readStack_entryFifoId_T_251 = _readStack_entryFifoId_T_243 + _readStack_entryFifoId_T_249; // @[ReadStack.scala 135:45]
  wire [4:0] _readStack_entryFifoId_T_253 = _readStack_entryFifoId_T_237 + _readStack_entryFifoId_T_251; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_255 = _axireqArb_io_in_16_valid_T_1 + _axireqArb_io_in_17_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_257 = _axireqArb_io_in_18_valid_T_1 + _axireqArb_io_in_19_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_259 = _readStack_entryFifoId_T_255 + _readStack_entryFifoId_T_257; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_261 = _axireqArb_io_in_20_valid_T_1 + _axireqArb_io_in_21_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_263 = _axireqArb_io_in_22_valid_T_1 + _axireqArb_io_in_23_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_265 = _readStack_entryFifoId_T_261 + _readStack_entryFifoId_T_263; // @[ReadStack.scala 135:45]
  wire [3:0] _readStack_entryFifoId_T_267 = _readStack_entryFifoId_T_259 + _readStack_entryFifoId_T_265; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_269 = _axireqArb_io_in_24_valid_T_1 + _axireqArb_io_in_25_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_271 = _axireqArb_io_in_26_valid_T_1 + _axireqArb_io_in_27_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_273 = _readStack_entryFifoId_T_269 + _readStack_entryFifoId_T_271; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_275 = _axireqArb_io_in_28_valid_T_1 + _axireqArb_io_in_29_valid_T_1; // @[ReadStack.scala 135:45]
  wire [1:0] _readStack_entryFifoId_T_277 = _axireqArb_io_in_30_valid_T_1 + _axireqArb_io_in_31_valid_T_1; // @[ReadStack.scala 135:45]
  wire [2:0] _readStack_entryFifoId_T_279 = _readStack_entryFifoId_T_275 + _readStack_entryFifoId_T_277; // @[ReadStack.scala 135:45]
  wire [3:0] _readStack_entryFifoId_T_281 = _readStack_entryFifoId_T_273 + _readStack_entryFifoId_T_279; // @[ReadStack.scala 135:45]
  wire [4:0] _readStack_entryFifoId_T_283 = _readStack_entryFifoId_T_267 + _readStack_entryFifoId_T_281; // @[ReadStack.scala 135:45]
  wire [5:0] _readStack_entryFifoId_T_285 = _readStack_entryFifoId_T_253 + _readStack_entryFifoId_T_283; // @[ReadStack.scala 135:45]
  wire [5:0] _GEN_416 = 5'h0 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_0_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_417 = 5'h1 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_1_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_418 = 5'h2 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_2_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_419 = 5'h3 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_3_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_420 = 5'h4 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_4_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_421 = 5'h5 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_5_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_422 = 5'h6 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_6_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_423 = 5'h7 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_7_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_424 = 5'h8 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_8_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_425 = 5'h9 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_9_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_426 = 5'ha == idxInsert ? _readStack_entryFifoId_T_285 : readStack_10_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_427 = 5'hb == idxInsert ? _readStack_entryFifoId_T_285 : readStack_11_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_428 = 5'hc == idxInsert ? _readStack_entryFifoId_T_285 : readStack_12_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_429 = 5'hd == idxInsert ? _readStack_entryFifoId_T_285 : readStack_13_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_430 = 5'he == idxInsert ? _readStack_entryFifoId_T_285 : readStack_14_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_431 = 5'hf == idxInsert ? _readStack_entryFifoId_T_285 : readStack_15_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_432 = 5'h10 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_16_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_433 = 5'h11 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_17_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_434 = 5'h12 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_18_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_435 = 5'h13 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_19_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_436 = 5'h14 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_20_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_437 = 5'h15 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_21_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_438 = 5'h16 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_22_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_439 = 5'h17 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_23_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_440 = 5'h18 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_24_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_441 = 5'h19 == idxInsert ? _readStack_entryFifoId_T_285 : readStack_25_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_442 = 5'h1a == idxInsert ? _readStack_entryFifoId_T_285 : readStack_26_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_443 = 5'h1b == idxInsert ? _readStack_entryFifoId_T_285 : readStack_27_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_444 = 5'h1c == idxInsert ? _readStack_entryFifoId_T_285 : readStack_28_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_445 = 5'h1d == idxInsert ? _readStack_entryFifoId_T_285 : readStack_29_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_446 = 5'h1e == idxInsert ? _readStack_entryFifoId_T_285 : readStack_30_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_447 = 5'h1f == idxInsert ? _readStack_entryFifoId_T_285 : readStack_31_entryFifoId; // @[ReadStack.scala 135:{27,27} 63:26]
  wire [5:0] _GEN_448 = _T_6 ? _GEN_416 : readStack_0_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_449 = _T_6 ? _GEN_417 : readStack_1_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_450 = _T_6 ? _GEN_418 : readStack_2_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_451 = _T_6 ? _GEN_419 : readStack_3_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_452 = _T_6 ? _GEN_420 : readStack_4_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_453 = _T_6 ? _GEN_421 : readStack_5_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_454 = _T_6 ? _GEN_422 : readStack_6_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_455 = _T_6 ? _GEN_423 : readStack_7_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_456 = _T_6 ? _GEN_424 : readStack_8_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_457 = _T_6 ? _GEN_425 : readStack_9_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_458 = _T_6 ? _GEN_426 : readStack_10_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_459 = _T_6 ? _GEN_427 : readStack_11_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_460 = _T_6 ? _GEN_428 : readStack_12_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_461 = _T_6 ? _GEN_429 : readStack_13_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_462 = _T_6 ? _GEN_430 : readStack_14_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_463 = _T_6 ? _GEN_431 : readStack_15_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_464 = _T_6 ? _GEN_432 : readStack_16_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_465 = _T_6 ? _GEN_433 : readStack_17_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_466 = _T_6 ? _GEN_434 : readStack_18_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_467 = _T_6 ? _GEN_435 : readStack_19_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_468 = _T_6 ? _GEN_436 : readStack_20_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_469 = _T_6 ? _GEN_437 : readStack_21_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_470 = _T_6 ? _GEN_438 : readStack_22_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_471 = _T_6 ? _GEN_439 : readStack_23_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_472 = _T_6 ? _GEN_440 : readStack_24_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_473 = _T_6 ? _GEN_441 : readStack_25_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_474 = _T_6 ? _GEN_442 : readStack_26_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_475 = _T_6 ? _GEN_443 : readStack_27_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_476 = _T_6 ? _GEN_444 : readStack_28_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_477 = _T_6 ? _GEN_445 : readStack_29_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_478 = _T_6 ? _GEN_446 : readStack_30_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_479 = _T_6 ? _GEN_447 : readStack_31_entryFifoId; // @[ReadStack.scala 132:5 63:26]
  wire [5:0] _GEN_480 = _T_2 ? _GEN_384 : _GEN_448; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_481 = _T_2 ? _GEN_385 : _GEN_449; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_482 = _T_2 ? _GEN_386 : _GEN_450; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_483 = _T_2 ? _GEN_387 : _GEN_451; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_484 = _T_2 ? _GEN_388 : _GEN_452; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_485 = _T_2 ? _GEN_389 : _GEN_453; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_486 = _T_2 ? _GEN_390 : _GEN_454; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_487 = _T_2 ? _GEN_391 : _GEN_455; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_488 = _T_2 ? _GEN_392 : _GEN_456; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_489 = _T_2 ? _GEN_393 : _GEN_457; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_490 = _T_2 ? _GEN_394 : _GEN_458; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_491 = _T_2 ? _GEN_395 : _GEN_459; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_492 = _T_2 ? _GEN_396 : _GEN_460; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_493 = _T_2 ? _GEN_397 : _GEN_461; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_494 = _T_2 ? _GEN_398 : _GEN_462; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_495 = _T_2 ? _GEN_399 : _GEN_463; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_496 = _T_2 ? _GEN_400 : _GEN_464; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_497 = _T_2 ? _GEN_401 : _GEN_465; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_498 = _T_2 ? _GEN_402 : _GEN_466; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_499 = _T_2 ? _GEN_403 : _GEN_467; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_500 = _T_2 ? _GEN_404 : _GEN_468; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_501 = _T_2 ? _GEN_405 : _GEN_469; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_502 = _T_2 ? _GEN_406 : _GEN_470; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_503 = _T_2 ? _GEN_407 : _GEN_471; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_504 = _T_2 ? _GEN_408 : _GEN_472; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_505 = _T_2 ? _GEN_409 : _GEN_473; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_506 = _T_2 ? _GEN_410 : _GEN_474; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_507 = _T_2 ? _GEN_411 : _GEN_475; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_508 = _T_2 ? _GEN_412 : _GEN_476; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_509 = _T_2 ? _GEN_413 : _GEN_477; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_510 = _T_2 ? _GEN_414 : _GEN_478; // @[ReadStack.scala 127:5]
  wire [5:0] _GEN_511 = _T_2 ? _GEN_415 : _GEN_479; // @[ReadStack.scala 127:5]
  wire [5:0] _readStack_0_entryFifoId_T_1 = readStack_0_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_1_entryFifoId_T_1 = readStack_1_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_2_entryFifoId_T_1 = readStack_2_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_3_entryFifoId_T_1 = readStack_3_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_4_entryFifoId_T_1 = readStack_4_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_5_entryFifoId_T_1 = readStack_5_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_6_entryFifoId_T_1 = readStack_6_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_7_entryFifoId_T_1 = readStack_7_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_8_entryFifoId_T_1 = readStack_8_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_9_entryFifoId_T_1 = readStack_9_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_10_entryFifoId_T_1 = readStack_10_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_11_entryFifoId_T_1 = readStack_11_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_12_entryFifoId_T_1 = readStack_12_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_13_entryFifoId_T_1 = readStack_13_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_14_entryFifoId_T_1 = readStack_14_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_15_entryFifoId_T_1 = readStack_15_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_16_entryFifoId_T_1 = readStack_16_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_17_entryFifoId_T_1 = readStack_17_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_18_entryFifoId_T_1 = readStack_18_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_19_entryFifoId_T_1 = readStack_19_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_20_entryFifoId_T_1 = readStack_20_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_21_entryFifoId_T_1 = readStack_21_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_22_entryFifoId_T_1 = readStack_22_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_23_entryFifoId_T_1 = readStack_23_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_24_entryFifoId_T_1 = readStack_24_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_25_entryFifoId_T_1 = readStack_25_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_26_entryFifoId_T_1 = readStack_26_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_27_entryFifoId_T_1 = readStack_27_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_28_entryFifoId_T_1 = readStack_28_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_29_entryFifoId_T_1 = readStack_29_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_30_entryFifoId_T_1 = readStack_30_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire [5:0] _readStack_31_entryFifoId_T_1 = readStack_31_entryFifoId - 6'h1; // @[ReadStack.scala 144:40]
  wire  _canReceive_T_1 = readStack_0_rvalid & _GEN_1184 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_3 = readStack_1_rvalid & _GEN_1185 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_5 = readStack_2_rvalid & _GEN_1186 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_7 = readStack_3_rvalid & _GEN_1187 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_9 = readStack_4_rvalid & _GEN_1188 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_11 = readStack_5_rvalid & _GEN_1189 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_13 = readStack_6_rvalid & _GEN_1190 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_15 = readStack_7_rvalid & _GEN_1191 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_17 = readStack_8_rvalid & _GEN_1192 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_19 = readStack_9_rvalid & _GEN_1193 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_21 = readStack_10_rvalid & _GEN_1194 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_23 = readStack_11_rvalid & _GEN_1195 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_25 = readStack_12_rvalid & _GEN_1196 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_27 = readStack_13_rvalid & _GEN_1197 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_29 = readStack_14_rvalid & _GEN_1198 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_31 = readStack_15_rvalid & _GEN_1199 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_33 = readStack_16_rvalid & _GEN_1200 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_35 = readStack_17_rvalid & _GEN_1201 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_37 = readStack_18_rvalid & _GEN_1202 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_39 = readStack_19_rvalid & _GEN_1203 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_41 = readStack_20_rvalid & _GEN_1204 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_43 = readStack_21_rvalid & _GEN_1205 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_45 = readStack_22_rvalid & _GEN_1206 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_47 = readStack_23_rvalid & _GEN_1207 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_49 = readStack_24_rvalid & _GEN_1208 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_51 = readStack_25_rvalid & _GEN_1209 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_53 = readStack_26_rvalid & _GEN_1210 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_55 = readStack_27_rvalid & _GEN_1211 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_57 = readStack_28_rvalid & _GEN_1212 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_59 = readStack_29_rvalid & _GEN_1213 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_61 = readStack_30_rvalid & _GEN_1214 == 3'h2; // @[ReadStack.scala 150:51]
  wire  _canReceive_T_63 = readStack_31_rvalid & _GEN_1215 == 3'h2; // @[ReadStack.scala 150:51]
  wire [7:0] canReceive_lo_lo = {_canReceive_T_49,_canReceive_T_51,_canReceive_T_53,_canReceive_T_55,_canReceive_T_57,
    _canReceive_T_59,_canReceive_T_61,_canReceive_T_63}; // @[Cat.scala 31:58]
  wire [15:0] canReceive_lo = {_canReceive_T_33,_canReceive_T_35,_canReceive_T_37,_canReceive_T_39,_canReceive_T_41,
    _canReceive_T_43,_canReceive_T_45,_canReceive_T_47,canReceive_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] canReceive_hi_lo = {_canReceive_T_17,_canReceive_T_19,_canReceive_T_21,_canReceive_T_23,_canReceive_T_25,
    _canReceive_T_27,_canReceive_T_29,_canReceive_T_31}; // @[Cat.scala 31:58]
  wire [31:0] _canReceive_T_64 = {_canReceive_T_1,_canReceive_T_3,_canReceive_T_5,_canReceive_T_7,_canReceive_T_9,
    _canReceive_T_11,_canReceive_T_13,_canReceive_T_15,canReceive_hi_lo,canReceive_lo}; // @[Cat.scala 31:58]
  wire [4:0] respEntryId = io_tlResp_in_d_bits_source[18:14]; // @[ReadStack.scala 153:29]
  wire  _readStack_respStatus_T = ~io_tlResp_in_d_bits_denied; // @[ReadStack.scala 157:27]
  wire [3:0] _readStack_respEntryId_respStatus = {{3'd0}, _readStack_respStatus_T}; // @[ReadStack.scala 157:{24,24}]
  wire  _T_72 = io_axiResp_out_r_ready & io_axiResp_out_r_valid; // @[Decoupled.scala 50:35]
  wire  _T_73 = alloc & _T_72; // @[ReadStack.scala 182:15]
  wire  _readStack_BeatFifoId_T_1 = readStack_0_rvalid & readStack_0_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_3 = readStack_1_rvalid & readStack_1_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_5 = readStack_2_rvalid & readStack_2_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_7 = readStack_3_rvalid & readStack_3_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_9 = readStack_4_rvalid & readStack_4_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_11 = readStack_5_rvalid & readStack_5_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_13 = readStack_6_rvalid & readStack_6_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_15 = readStack_7_rvalid & readStack_7_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_17 = readStack_8_rvalid & readStack_8_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_19 = readStack_9_rvalid & readStack_9_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_21 = readStack_10_rvalid & readStack_10_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_23 = readStack_11_rvalid & readStack_11_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_25 = readStack_12_rvalid & readStack_12_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_27 = readStack_13_rvalid & readStack_13_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_29 = readStack_14_rvalid & readStack_14_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_31 = readStack_15_rvalid & readStack_15_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_33 = readStack_16_rvalid & readStack_16_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_35 = readStack_17_rvalid & readStack_17_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_37 = readStack_18_rvalid & readStack_18_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_39 = readStack_19_rvalid & readStack_19_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_41 = readStack_20_rvalid & readStack_20_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_43 = readStack_21_rvalid & readStack_21_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_45 = readStack_22_rvalid & readStack_22_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_47 = readStack_23_rvalid & readStack_23_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_49 = readStack_24_rvalid & readStack_24_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_51 = readStack_25_rvalid & readStack_25_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_53 = readStack_26_rvalid & readStack_26_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_55 = readStack_27_rvalid & readStack_27_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_57 = readStack_28_rvalid & readStack_28_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_59 = readStack_29_rvalid & readStack_29_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_61 = readStack_30_rvalid & readStack_30_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire  _readStack_BeatFifoId_T_63 = readStack_31_rvalid & readStack_31_arid == io_axiReq_in_ar_bits_id; // @[ReadStack.scala 185:70]
  wire [7:0] readStack_BeatFifoId_lo_lo = {_readStack_BeatFifoId_T_49,_readStack_BeatFifoId_T_51,
    _readStack_BeatFifoId_T_53,_readStack_BeatFifoId_T_55,_readStack_BeatFifoId_T_57,_readStack_BeatFifoId_T_59,
    _readStack_BeatFifoId_T_61,_readStack_BeatFifoId_T_63}; // @[Cat.scala 31:58]
  wire [15:0] readStack_BeatFifoId_lo = {_readStack_BeatFifoId_T_33,_readStack_BeatFifoId_T_35,
    _readStack_BeatFifoId_T_37,_readStack_BeatFifoId_T_39,_readStack_BeatFifoId_T_41,_readStack_BeatFifoId_T_43,
    _readStack_BeatFifoId_T_45,_readStack_BeatFifoId_T_47,readStack_BeatFifoId_lo_lo}; // @[Cat.scala 31:58]
  wire [7:0] readStack_BeatFifoId_hi_lo = {_readStack_BeatFifoId_T_17,_readStack_BeatFifoId_T_19,
    _readStack_BeatFifoId_T_21,_readStack_BeatFifoId_T_23,_readStack_BeatFifoId_T_25,_readStack_BeatFifoId_T_27,
    _readStack_BeatFifoId_T_29,_readStack_BeatFifoId_T_31}; // @[Cat.scala 31:58]
  wire [31:0] _readStack_BeatFifoId_T_64 = {_readStack_BeatFifoId_T_1,_readStack_BeatFifoId_T_3,
    _readStack_BeatFifoId_T_5,_readStack_BeatFifoId_T_7,_readStack_BeatFifoId_T_9,_readStack_BeatFifoId_T_11,
    _readStack_BeatFifoId_T_13,_readStack_BeatFifoId_T_15,readStack_BeatFifoId_hi_lo,readStack_BeatFifoId_lo}; // @[Cat.scala 31:58]
  wire [1:0] _readStack_BeatFifoId_T_97 = _readStack_BeatFifoId_T_64[0] + _readStack_BeatFifoId_T_64[1]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_99 = _readStack_BeatFifoId_T_64[2] + _readStack_BeatFifoId_T_64[3]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_101 = _readStack_BeatFifoId_T_97 + _readStack_BeatFifoId_T_99; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_103 = _readStack_BeatFifoId_T_64[4] + _readStack_BeatFifoId_T_64[5]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_105 = _readStack_BeatFifoId_T_64[6] + _readStack_BeatFifoId_T_64[7]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_107 = _readStack_BeatFifoId_T_103 + _readStack_BeatFifoId_T_105; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_BeatFifoId_T_109 = _readStack_BeatFifoId_T_101 + _readStack_BeatFifoId_T_107; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_111 = _readStack_BeatFifoId_T_64[8] + _readStack_BeatFifoId_T_64[9]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_113 = _readStack_BeatFifoId_T_64[10] + _readStack_BeatFifoId_T_64[11]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_115 = _readStack_BeatFifoId_T_111 + _readStack_BeatFifoId_T_113; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_117 = _readStack_BeatFifoId_T_64[12] + _readStack_BeatFifoId_T_64[13]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_119 = _readStack_BeatFifoId_T_64[14] + _readStack_BeatFifoId_T_64[15]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_121 = _readStack_BeatFifoId_T_117 + _readStack_BeatFifoId_T_119; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_BeatFifoId_T_123 = _readStack_BeatFifoId_T_115 + _readStack_BeatFifoId_T_121; // @[Bitwise.scala 48:55]
  wire [4:0] _readStack_BeatFifoId_T_125 = _readStack_BeatFifoId_T_109 + _readStack_BeatFifoId_T_123; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_127 = _readStack_BeatFifoId_T_64[16] + _readStack_BeatFifoId_T_64[17]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_129 = _readStack_BeatFifoId_T_64[18] + _readStack_BeatFifoId_T_64[19]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_131 = _readStack_BeatFifoId_T_127 + _readStack_BeatFifoId_T_129; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_133 = _readStack_BeatFifoId_T_64[20] + _readStack_BeatFifoId_T_64[21]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_135 = _readStack_BeatFifoId_T_64[22] + _readStack_BeatFifoId_T_64[23]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_137 = _readStack_BeatFifoId_T_133 + _readStack_BeatFifoId_T_135; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_BeatFifoId_T_139 = _readStack_BeatFifoId_T_131 + _readStack_BeatFifoId_T_137; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_141 = _readStack_BeatFifoId_T_64[24] + _readStack_BeatFifoId_T_64[25]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_143 = _readStack_BeatFifoId_T_64[26] + _readStack_BeatFifoId_T_64[27]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_145 = _readStack_BeatFifoId_T_141 + _readStack_BeatFifoId_T_143; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_147 = _readStack_BeatFifoId_T_64[28] + _readStack_BeatFifoId_T_64[29]; // @[Bitwise.scala 48:55]
  wire [1:0] _readStack_BeatFifoId_T_149 = _readStack_BeatFifoId_T_64[30] + _readStack_BeatFifoId_T_64[31]; // @[Bitwise.scala 48:55]
  wire [2:0] _readStack_BeatFifoId_T_151 = _readStack_BeatFifoId_T_147 + _readStack_BeatFifoId_T_149; // @[Bitwise.scala 48:55]
  wire [3:0] _readStack_BeatFifoId_T_153 = _readStack_BeatFifoId_T_145 + _readStack_BeatFifoId_T_151; // @[Bitwise.scala 48:55]
  wire [4:0] _readStack_BeatFifoId_T_155 = _readStack_BeatFifoId_T_139 + _readStack_BeatFifoId_T_153; // @[Bitwise.scala 48:55]
  wire [5:0] _readStack_BeatFifoId_T_157 = _readStack_BeatFifoId_T_125 + _readStack_BeatFifoId_T_155; // @[Bitwise.scala 48:55]
  wire [5:0] _readStack_BeatFifoId_T_160 = _readStack_BeatFifoId_T_157 - 6'h1; // @[ReadStack.scala 185:113]
  wire [5:0] _GEN_800 = 5'h0 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_0_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_801 = 5'h1 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_1_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_802 = 5'h2 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_2_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_803 = 5'h3 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_3_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_804 = 5'h4 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_4_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_805 = 5'h5 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_5_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_806 = 5'h6 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_6_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_807 = 5'h7 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_7_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_808 = 5'h8 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_8_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_809 = 5'h9 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_9_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_810 = 5'ha == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_10_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_811 = 5'hb == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_11_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_812 = 5'hc == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_12_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_813 = 5'hd == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_13_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_814 = 5'he == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_14_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_815 = 5'hf == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_15_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_816 = 5'h10 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_16_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_817 = 5'h11 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_17_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_818 = 5'h12 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_18_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_819 = 5'h13 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_19_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_820 = 5'h14 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_20_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_821 = 5'h15 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_21_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_822 = 5'h16 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_22_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_823 = 5'h17 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_23_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_824 = 5'h18 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_24_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_825 = 5'h19 == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_25_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_826 = 5'h1a == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_26_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_827 = 5'h1b == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_27_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_828 = 5'h1c == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_28_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_829 = 5'h1d == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_29_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_830 = 5'h1e == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_30_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire [5:0] _GEN_831 = 5'h1f == idxInsert ? _readStack_BeatFifoId_T_160 : readStack_31_BeatFifoId; // @[ReadStack.scala 185:{26,26} 63:26]
  wire  _T_76 = alloc & ~_T_72; // @[ReadStack.scala 186:25]
  wire [1:0] _readStack_BeatFifoId_T_225 = _readStack_BeatFifoId_T_1 + _readStack_BeatFifoId_T_3; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_227 = _readStack_BeatFifoId_T_5 + _readStack_BeatFifoId_T_7; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_229 = _readStack_BeatFifoId_T_225 + _readStack_BeatFifoId_T_227; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_231 = _readStack_BeatFifoId_T_9 + _readStack_BeatFifoId_T_11; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_233 = _readStack_BeatFifoId_T_13 + _readStack_BeatFifoId_T_15; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_235 = _readStack_BeatFifoId_T_231 + _readStack_BeatFifoId_T_233; // @[ReadStack.scala 189:46]
  wire [3:0] _readStack_BeatFifoId_T_237 = _readStack_BeatFifoId_T_229 + _readStack_BeatFifoId_T_235; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_239 = _readStack_BeatFifoId_T_17 + _readStack_BeatFifoId_T_19; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_241 = _readStack_BeatFifoId_T_21 + _readStack_BeatFifoId_T_23; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_243 = _readStack_BeatFifoId_T_239 + _readStack_BeatFifoId_T_241; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_245 = _readStack_BeatFifoId_T_25 + _readStack_BeatFifoId_T_27; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_247 = _readStack_BeatFifoId_T_29 + _readStack_BeatFifoId_T_31; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_249 = _readStack_BeatFifoId_T_245 + _readStack_BeatFifoId_T_247; // @[ReadStack.scala 189:46]
  wire [3:0] _readStack_BeatFifoId_T_251 = _readStack_BeatFifoId_T_243 + _readStack_BeatFifoId_T_249; // @[ReadStack.scala 189:46]
  wire [4:0] _readStack_BeatFifoId_T_253 = _readStack_BeatFifoId_T_237 + _readStack_BeatFifoId_T_251; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_255 = _readStack_BeatFifoId_T_33 + _readStack_BeatFifoId_T_35; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_257 = _readStack_BeatFifoId_T_37 + _readStack_BeatFifoId_T_39; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_259 = _readStack_BeatFifoId_T_255 + _readStack_BeatFifoId_T_257; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_261 = _readStack_BeatFifoId_T_41 + _readStack_BeatFifoId_T_43; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_263 = _readStack_BeatFifoId_T_45 + _readStack_BeatFifoId_T_47; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_265 = _readStack_BeatFifoId_T_261 + _readStack_BeatFifoId_T_263; // @[ReadStack.scala 189:46]
  wire [3:0] _readStack_BeatFifoId_T_267 = _readStack_BeatFifoId_T_259 + _readStack_BeatFifoId_T_265; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_269 = _readStack_BeatFifoId_T_49 + _readStack_BeatFifoId_T_51; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_271 = _readStack_BeatFifoId_T_53 + _readStack_BeatFifoId_T_55; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_273 = _readStack_BeatFifoId_T_269 + _readStack_BeatFifoId_T_271; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_275 = _readStack_BeatFifoId_T_57 + _readStack_BeatFifoId_T_59; // @[ReadStack.scala 189:46]
  wire [1:0] _readStack_BeatFifoId_T_277 = _readStack_BeatFifoId_T_61 + _readStack_BeatFifoId_T_63; // @[ReadStack.scala 189:46]
  wire [2:0] _readStack_BeatFifoId_T_279 = _readStack_BeatFifoId_T_275 + _readStack_BeatFifoId_T_277; // @[ReadStack.scala 189:46]
  wire [3:0] _readStack_BeatFifoId_T_281 = _readStack_BeatFifoId_T_273 + _readStack_BeatFifoId_T_279; // @[ReadStack.scala 189:46]
  wire [4:0] _readStack_BeatFifoId_T_283 = _readStack_BeatFifoId_T_267 + _readStack_BeatFifoId_T_281; // @[ReadStack.scala 189:46]
  wire [5:0] _readStack_BeatFifoId_T_285 = _readStack_BeatFifoId_T_253 + _readStack_BeatFifoId_T_283; // @[ReadStack.scala 189:46]
  wire [5:0] _GEN_832 = 5'h0 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_0_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_833 = 5'h1 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_1_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_834 = 5'h2 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_2_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_835 = 5'h3 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_3_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_836 = 5'h4 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_4_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_837 = 5'h5 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_5_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_838 = 5'h6 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_6_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_839 = 5'h7 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_7_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_840 = 5'h8 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_8_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_841 = 5'h9 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_9_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_842 = 5'ha == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_10_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_843 = 5'hb == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_11_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_844 = 5'hc == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_12_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_845 = 5'hd == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_13_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_846 = 5'he == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_14_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_847 = 5'hf == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_15_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_848 = 5'h10 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_16_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_849 = 5'h11 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_17_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_850 = 5'h12 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_18_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_851 = 5'h13 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_19_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_852 = 5'h14 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_20_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_853 = 5'h15 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_21_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_854 = 5'h16 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_22_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_855 = 5'h17 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_23_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_856 = 5'h18 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_24_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_857 = 5'h19 == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_25_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_858 = 5'h1a == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_26_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_859 = 5'h1b == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_27_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_860 = 5'h1c == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_28_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_861 = 5'h1d == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_29_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_862 = 5'h1e == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_30_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_863 = 5'h1f == idxInsert ? _readStack_BeatFifoId_T_285 : readStack_31_BeatFifoId; // @[ReadStack.scala 189:{28,28} 63:26]
  wire [5:0] _GEN_864 = _T_76 ? _GEN_832 : readStack_0_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_865 = _T_76 ? _GEN_833 : readStack_1_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_866 = _T_76 ? _GEN_834 : readStack_2_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_867 = _T_76 ? _GEN_835 : readStack_3_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_868 = _T_76 ? _GEN_836 : readStack_4_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_869 = _T_76 ? _GEN_837 : readStack_5_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_870 = _T_76 ? _GEN_838 : readStack_6_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_871 = _T_76 ? _GEN_839 : readStack_7_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_872 = _T_76 ? _GEN_840 : readStack_8_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_873 = _T_76 ? _GEN_841 : readStack_9_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_874 = _T_76 ? _GEN_842 : readStack_10_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_875 = _T_76 ? _GEN_843 : readStack_11_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_876 = _T_76 ? _GEN_844 : readStack_12_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_877 = _T_76 ? _GEN_845 : readStack_13_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_878 = _T_76 ? _GEN_846 : readStack_14_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_879 = _T_76 ? _GEN_847 : readStack_15_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_880 = _T_76 ? _GEN_848 : readStack_16_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_881 = _T_76 ? _GEN_849 : readStack_17_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_882 = _T_76 ? _GEN_850 : readStack_18_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_883 = _T_76 ? _GEN_851 : readStack_19_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_884 = _T_76 ? _GEN_852 : readStack_20_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_885 = _T_76 ? _GEN_853 : readStack_21_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_886 = _T_76 ? _GEN_854 : readStack_22_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_887 = _T_76 ? _GEN_855 : readStack_23_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_888 = _T_76 ? _GEN_856 : readStack_24_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_889 = _T_76 ? _GEN_857 : readStack_25_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_890 = _T_76 ? _GEN_858 : readStack_26_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_891 = _T_76 ? _GEN_859 : readStack_27_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_892 = _T_76 ? _GEN_860 : readStack_28_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_893 = _T_76 ? _GEN_861 : readStack_29_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_894 = _T_76 ? _GEN_862 : readStack_30_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_895 = _T_76 ? _GEN_863 : readStack_31_BeatFifoId; // @[ReadStack.scala 187:9 63:26]
  wire [5:0] _GEN_896 = _T_73 ? _GEN_800 : _GEN_864; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_897 = _T_73 ? _GEN_801 : _GEN_865; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_898 = _T_73 ? _GEN_802 : _GEN_866; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_899 = _T_73 ? _GEN_803 : _GEN_867; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_900 = _T_73 ? _GEN_804 : _GEN_868; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_901 = _T_73 ? _GEN_805 : _GEN_869; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_902 = _T_73 ? _GEN_806 : _GEN_870; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_903 = _T_73 ? _GEN_807 : _GEN_871; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_904 = _T_73 ? _GEN_808 : _GEN_872; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_905 = _T_73 ? _GEN_809 : _GEN_873; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_906 = _T_73 ? _GEN_810 : _GEN_874; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_907 = _T_73 ? _GEN_811 : _GEN_875; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_908 = _T_73 ? _GEN_812 : _GEN_876; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_909 = _T_73 ? _GEN_813 : _GEN_877; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_910 = _T_73 ? _GEN_814 : _GEN_878; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_911 = _T_73 ? _GEN_815 : _GEN_879; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_912 = _T_73 ? _GEN_816 : _GEN_880; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_913 = _T_73 ? _GEN_817 : _GEN_881; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_914 = _T_73 ? _GEN_818 : _GEN_882; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_915 = _T_73 ? _GEN_819 : _GEN_883; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_916 = _T_73 ? _GEN_820 : _GEN_884; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_917 = _T_73 ? _GEN_821 : _GEN_885; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_918 = _T_73 ? _GEN_822 : _GEN_886; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_919 = _T_73 ? _GEN_823 : _GEN_887; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_920 = _T_73 ? _GEN_824 : _GEN_888; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_921 = _T_73 ? _GEN_825 : _GEN_889; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_922 = _T_73 ? _GEN_826 : _GEN_890; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_923 = _T_73 ? _GEN_827 : _GEN_891; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_924 = _T_73 ? _GEN_828 : _GEN_892; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_925 = _T_73 ? _GEN_829 : _GEN_893; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_926 = _T_73 ? _GEN_830 : _GEN_894; // @[ReadStack.scala 183:7]
  wire [5:0] _GEN_927 = _T_73 ? _GEN_831 : _GEN_895; // @[ReadStack.scala 183:7]
  wire [13:0] _GEN_993 = 5'h1 == axirespArb_io_chosen ? readStack_1_arid : readStack_0_arid; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_994 = 5'h2 == axirespArb_io_chosen ? readStack_2_arid : _GEN_993; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_995 = 5'h3 == axirespArb_io_chosen ? readStack_3_arid : _GEN_994; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_996 = 5'h4 == axirespArb_io_chosen ? readStack_4_arid : _GEN_995; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_997 = 5'h5 == axirespArb_io_chosen ? readStack_5_arid : _GEN_996; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_998 = 5'h6 == axirespArb_io_chosen ? readStack_6_arid : _GEN_997; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_999 = 5'h7 == axirespArb_io_chosen ? readStack_7_arid : _GEN_998; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1000 = 5'h8 == axirespArb_io_chosen ? readStack_8_arid : _GEN_999; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1001 = 5'h9 == axirespArb_io_chosen ? readStack_9_arid : _GEN_1000; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1002 = 5'ha == axirespArb_io_chosen ? readStack_10_arid : _GEN_1001; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1003 = 5'hb == axirespArb_io_chosen ? readStack_11_arid : _GEN_1002; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1004 = 5'hc == axirespArb_io_chosen ? readStack_12_arid : _GEN_1003; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1005 = 5'hd == axirespArb_io_chosen ? readStack_13_arid : _GEN_1004; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1006 = 5'he == axirespArb_io_chosen ? readStack_14_arid : _GEN_1005; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1007 = 5'hf == axirespArb_io_chosen ? readStack_15_arid : _GEN_1006; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1008 = 5'h10 == axirespArb_io_chosen ? readStack_16_arid : _GEN_1007; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1009 = 5'h11 == axirespArb_io_chosen ? readStack_17_arid : _GEN_1008; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1010 = 5'h12 == axirespArb_io_chosen ? readStack_18_arid : _GEN_1009; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1011 = 5'h13 == axirespArb_io_chosen ? readStack_19_arid : _GEN_1010; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1012 = 5'h14 == axirespArb_io_chosen ? readStack_20_arid : _GEN_1011; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1013 = 5'h15 == axirespArb_io_chosen ? readStack_21_arid : _GEN_1012; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1014 = 5'h16 == axirespArb_io_chosen ? readStack_22_arid : _GEN_1013; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1015 = 5'h17 == axirespArb_io_chosen ? readStack_23_arid : _GEN_1014; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1016 = 5'h18 == axirespArb_io_chosen ? readStack_24_arid : _GEN_1015; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1017 = 5'h19 == axirespArb_io_chosen ? readStack_25_arid : _GEN_1016; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1018 = 5'h1a == axirespArb_io_chosen ? readStack_26_arid : _GEN_1017; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1019 = 5'h1b == axirespArb_io_chosen ? readStack_27_arid : _GEN_1018; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1020 = 5'h1c == axirespArb_io_chosen ? readStack_28_arid : _GEN_1019; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1021 = 5'h1d == axirespArb_io_chosen ? readStack_29_arid : _GEN_1020; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1022 = 5'h1e == axirespArb_io_chosen ? readStack_30_arid : _GEN_1021; // @[ReadStack.scala 196:{35,35}]
  wire [13:0] _GEN_1023 = 5'h1f == axirespArb_io_chosen ? readStack_31_arid : _GEN_1022; // @[ReadStack.scala 196:{35,35}]
  wire [5:0] _readStack_0_BeatFifoId_T_1 = readStack_0_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_1_BeatFifoId_T_1 = readStack_1_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_2_BeatFifoId_T_1 = readStack_2_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_3_BeatFifoId_T_1 = readStack_3_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_4_BeatFifoId_T_1 = readStack_4_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_5_BeatFifoId_T_1 = readStack_5_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_6_BeatFifoId_T_1 = readStack_6_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_7_BeatFifoId_T_1 = readStack_7_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_8_BeatFifoId_T_1 = readStack_8_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_9_BeatFifoId_T_1 = readStack_9_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_10_BeatFifoId_T_1 = readStack_10_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_11_BeatFifoId_T_1 = readStack_11_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_12_BeatFifoId_T_1 = readStack_12_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_13_BeatFifoId_T_1 = readStack_13_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_14_BeatFifoId_T_1 = readStack_14_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_15_BeatFifoId_T_1 = readStack_15_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_16_BeatFifoId_T_1 = readStack_16_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_17_BeatFifoId_T_1 = readStack_17_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_18_BeatFifoId_T_1 = readStack_18_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_19_BeatFifoId_T_1 = readStack_19_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_20_BeatFifoId_T_1 = readStack_20_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_21_BeatFifoId_T_1 = readStack_21_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_22_BeatFifoId_T_1 = readStack_22_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_23_BeatFifoId_T_1 = readStack_23_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_24_BeatFifoId_T_1 = readStack_24_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_25_BeatFifoId_T_1 = readStack_25_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_26_BeatFifoId_T_1 = readStack_26_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_27_BeatFifoId_T_1 = readStack_27_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_28_BeatFifoId_T_1 = readStack_28_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_29_BeatFifoId_T_1 = readStack_29_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_30_BeatFifoId_T_1 = readStack_30_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  wire [5:0] _readStack_31_BeatFifoId_T_1 = readStack_31_BeatFifoId - 6'h1; // @[ReadStack.scala 197:42]
  Arbiter axireqArb ( // @[ReadStack.scala 65:25]
    .io_in_0_valid(axireqArb_io_in_0_valid),
    .io_in_0_bits_raddress(axireqArb_io_in_0_bits_raddress),
    .io_in_0_bits_entryid(axireqArb_io_in_0_bits_entryid),
    .io_in_0_bits_arid(axireqArb_io_in_0_bits_arid),
    .io_in_0_bits_ardata(axireqArb_io_in_0_bits_ardata),
    .io_in_0_bits_respStatus(axireqArb_io_in_0_bits_respStatus),
    .io_in_0_bits_rsize(axireqArb_io_in_0_bits_rsize),
    .io_in_1_valid(axireqArb_io_in_1_valid),
    .io_in_1_bits_raddress(axireqArb_io_in_1_bits_raddress),
    .io_in_1_bits_entryid(axireqArb_io_in_1_bits_entryid),
    .io_in_1_bits_arid(axireqArb_io_in_1_bits_arid),
    .io_in_1_bits_ardata(axireqArb_io_in_1_bits_ardata),
    .io_in_1_bits_respStatus(axireqArb_io_in_1_bits_respStatus),
    .io_in_1_bits_rsize(axireqArb_io_in_1_bits_rsize),
    .io_in_2_valid(axireqArb_io_in_2_valid),
    .io_in_2_bits_raddress(axireqArb_io_in_2_bits_raddress),
    .io_in_2_bits_entryid(axireqArb_io_in_2_bits_entryid),
    .io_in_2_bits_arid(axireqArb_io_in_2_bits_arid),
    .io_in_2_bits_ardata(axireqArb_io_in_2_bits_ardata),
    .io_in_2_bits_respStatus(axireqArb_io_in_2_bits_respStatus),
    .io_in_2_bits_rsize(axireqArb_io_in_2_bits_rsize),
    .io_in_3_valid(axireqArb_io_in_3_valid),
    .io_in_3_bits_raddress(axireqArb_io_in_3_bits_raddress),
    .io_in_3_bits_entryid(axireqArb_io_in_3_bits_entryid),
    .io_in_3_bits_arid(axireqArb_io_in_3_bits_arid),
    .io_in_3_bits_ardata(axireqArb_io_in_3_bits_ardata),
    .io_in_3_bits_respStatus(axireqArb_io_in_3_bits_respStatus),
    .io_in_3_bits_rsize(axireqArb_io_in_3_bits_rsize),
    .io_in_4_valid(axireqArb_io_in_4_valid),
    .io_in_4_bits_raddress(axireqArb_io_in_4_bits_raddress),
    .io_in_4_bits_entryid(axireqArb_io_in_4_bits_entryid),
    .io_in_4_bits_arid(axireqArb_io_in_4_bits_arid),
    .io_in_4_bits_ardata(axireqArb_io_in_4_bits_ardata),
    .io_in_4_bits_respStatus(axireqArb_io_in_4_bits_respStatus),
    .io_in_4_bits_rsize(axireqArb_io_in_4_bits_rsize),
    .io_in_5_valid(axireqArb_io_in_5_valid),
    .io_in_5_bits_raddress(axireqArb_io_in_5_bits_raddress),
    .io_in_5_bits_entryid(axireqArb_io_in_5_bits_entryid),
    .io_in_5_bits_arid(axireqArb_io_in_5_bits_arid),
    .io_in_5_bits_ardata(axireqArb_io_in_5_bits_ardata),
    .io_in_5_bits_respStatus(axireqArb_io_in_5_bits_respStatus),
    .io_in_5_bits_rsize(axireqArb_io_in_5_bits_rsize),
    .io_in_6_valid(axireqArb_io_in_6_valid),
    .io_in_6_bits_raddress(axireqArb_io_in_6_bits_raddress),
    .io_in_6_bits_entryid(axireqArb_io_in_6_bits_entryid),
    .io_in_6_bits_arid(axireqArb_io_in_6_bits_arid),
    .io_in_6_bits_ardata(axireqArb_io_in_6_bits_ardata),
    .io_in_6_bits_respStatus(axireqArb_io_in_6_bits_respStatus),
    .io_in_6_bits_rsize(axireqArb_io_in_6_bits_rsize),
    .io_in_7_valid(axireqArb_io_in_7_valid),
    .io_in_7_bits_raddress(axireqArb_io_in_7_bits_raddress),
    .io_in_7_bits_entryid(axireqArb_io_in_7_bits_entryid),
    .io_in_7_bits_arid(axireqArb_io_in_7_bits_arid),
    .io_in_7_bits_ardata(axireqArb_io_in_7_bits_ardata),
    .io_in_7_bits_respStatus(axireqArb_io_in_7_bits_respStatus),
    .io_in_7_bits_rsize(axireqArb_io_in_7_bits_rsize),
    .io_in_8_valid(axireqArb_io_in_8_valid),
    .io_in_8_bits_raddress(axireqArb_io_in_8_bits_raddress),
    .io_in_8_bits_entryid(axireqArb_io_in_8_bits_entryid),
    .io_in_8_bits_arid(axireqArb_io_in_8_bits_arid),
    .io_in_8_bits_ardata(axireqArb_io_in_8_bits_ardata),
    .io_in_8_bits_respStatus(axireqArb_io_in_8_bits_respStatus),
    .io_in_8_bits_rsize(axireqArb_io_in_8_bits_rsize),
    .io_in_9_valid(axireqArb_io_in_9_valid),
    .io_in_9_bits_raddress(axireqArb_io_in_9_bits_raddress),
    .io_in_9_bits_entryid(axireqArb_io_in_9_bits_entryid),
    .io_in_9_bits_arid(axireqArb_io_in_9_bits_arid),
    .io_in_9_bits_ardata(axireqArb_io_in_9_bits_ardata),
    .io_in_9_bits_respStatus(axireqArb_io_in_9_bits_respStatus),
    .io_in_9_bits_rsize(axireqArb_io_in_9_bits_rsize),
    .io_in_10_valid(axireqArb_io_in_10_valid),
    .io_in_10_bits_raddress(axireqArb_io_in_10_bits_raddress),
    .io_in_10_bits_entryid(axireqArb_io_in_10_bits_entryid),
    .io_in_10_bits_arid(axireqArb_io_in_10_bits_arid),
    .io_in_10_bits_ardata(axireqArb_io_in_10_bits_ardata),
    .io_in_10_bits_respStatus(axireqArb_io_in_10_bits_respStatus),
    .io_in_10_bits_rsize(axireqArb_io_in_10_bits_rsize),
    .io_in_11_valid(axireqArb_io_in_11_valid),
    .io_in_11_bits_raddress(axireqArb_io_in_11_bits_raddress),
    .io_in_11_bits_entryid(axireqArb_io_in_11_bits_entryid),
    .io_in_11_bits_arid(axireqArb_io_in_11_bits_arid),
    .io_in_11_bits_ardata(axireqArb_io_in_11_bits_ardata),
    .io_in_11_bits_respStatus(axireqArb_io_in_11_bits_respStatus),
    .io_in_11_bits_rsize(axireqArb_io_in_11_bits_rsize),
    .io_in_12_valid(axireqArb_io_in_12_valid),
    .io_in_12_bits_raddress(axireqArb_io_in_12_bits_raddress),
    .io_in_12_bits_entryid(axireqArb_io_in_12_bits_entryid),
    .io_in_12_bits_arid(axireqArb_io_in_12_bits_arid),
    .io_in_12_bits_ardata(axireqArb_io_in_12_bits_ardata),
    .io_in_12_bits_respStatus(axireqArb_io_in_12_bits_respStatus),
    .io_in_12_bits_rsize(axireqArb_io_in_12_bits_rsize),
    .io_in_13_valid(axireqArb_io_in_13_valid),
    .io_in_13_bits_raddress(axireqArb_io_in_13_bits_raddress),
    .io_in_13_bits_entryid(axireqArb_io_in_13_bits_entryid),
    .io_in_13_bits_arid(axireqArb_io_in_13_bits_arid),
    .io_in_13_bits_ardata(axireqArb_io_in_13_bits_ardata),
    .io_in_13_bits_respStatus(axireqArb_io_in_13_bits_respStatus),
    .io_in_13_bits_rsize(axireqArb_io_in_13_bits_rsize),
    .io_in_14_valid(axireqArb_io_in_14_valid),
    .io_in_14_bits_raddress(axireqArb_io_in_14_bits_raddress),
    .io_in_14_bits_entryid(axireqArb_io_in_14_bits_entryid),
    .io_in_14_bits_arid(axireqArb_io_in_14_bits_arid),
    .io_in_14_bits_ardata(axireqArb_io_in_14_bits_ardata),
    .io_in_14_bits_respStatus(axireqArb_io_in_14_bits_respStatus),
    .io_in_14_bits_rsize(axireqArb_io_in_14_bits_rsize),
    .io_in_15_valid(axireqArb_io_in_15_valid),
    .io_in_15_bits_raddress(axireqArb_io_in_15_bits_raddress),
    .io_in_15_bits_entryid(axireqArb_io_in_15_bits_entryid),
    .io_in_15_bits_arid(axireqArb_io_in_15_bits_arid),
    .io_in_15_bits_ardata(axireqArb_io_in_15_bits_ardata),
    .io_in_15_bits_respStatus(axireqArb_io_in_15_bits_respStatus),
    .io_in_15_bits_rsize(axireqArb_io_in_15_bits_rsize),
    .io_in_16_valid(axireqArb_io_in_16_valid),
    .io_in_16_bits_raddress(axireqArb_io_in_16_bits_raddress),
    .io_in_16_bits_entryid(axireqArb_io_in_16_bits_entryid),
    .io_in_16_bits_arid(axireqArb_io_in_16_bits_arid),
    .io_in_16_bits_ardata(axireqArb_io_in_16_bits_ardata),
    .io_in_16_bits_respStatus(axireqArb_io_in_16_bits_respStatus),
    .io_in_16_bits_rsize(axireqArb_io_in_16_bits_rsize),
    .io_in_17_valid(axireqArb_io_in_17_valid),
    .io_in_17_bits_raddress(axireqArb_io_in_17_bits_raddress),
    .io_in_17_bits_entryid(axireqArb_io_in_17_bits_entryid),
    .io_in_17_bits_arid(axireqArb_io_in_17_bits_arid),
    .io_in_17_bits_ardata(axireqArb_io_in_17_bits_ardata),
    .io_in_17_bits_respStatus(axireqArb_io_in_17_bits_respStatus),
    .io_in_17_bits_rsize(axireqArb_io_in_17_bits_rsize),
    .io_in_18_valid(axireqArb_io_in_18_valid),
    .io_in_18_bits_raddress(axireqArb_io_in_18_bits_raddress),
    .io_in_18_bits_entryid(axireqArb_io_in_18_bits_entryid),
    .io_in_18_bits_arid(axireqArb_io_in_18_bits_arid),
    .io_in_18_bits_ardata(axireqArb_io_in_18_bits_ardata),
    .io_in_18_bits_respStatus(axireqArb_io_in_18_bits_respStatus),
    .io_in_18_bits_rsize(axireqArb_io_in_18_bits_rsize),
    .io_in_19_valid(axireqArb_io_in_19_valid),
    .io_in_19_bits_raddress(axireqArb_io_in_19_bits_raddress),
    .io_in_19_bits_entryid(axireqArb_io_in_19_bits_entryid),
    .io_in_19_bits_arid(axireqArb_io_in_19_bits_arid),
    .io_in_19_bits_ardata(axireqArb_io_in_19_bits_ardata),
    .io_in_19_bits_respStatus(axireqArb_io_in_19_bits_respStatus),
    .io_in_19_bits_rsize(axireqArb_io_in_19_bits_rsize),
    .io_in_20_valid(axireqArb_io_in_20_valid),
    .io_in_20_bits_raddress(axireqArb_io_in_20_bits_raddress),
    .io_in_20_bits_entryid(axireqArb_io_in_20_bits_entryid),
    .io_in_20_bits_arid(axireqArb_io_in_20_bits_arid),
    .io_in_20_bits_ardata(axireqArb_io_in_20_bits_ardata),
    .io_in_20_bits_respStatus(axireqArb_io_in_20_bits_respStatus),
    .io_in_20_bits_rsize(axireqArb_io_in_20_bits_rsize),
    .io_in_21_valid(axireqArb_io_in_21_valid),
    .io_in_21_bits_raddress(axireqArb_io_in_21_bits_raddress),
    .io_in_21_bits_entryid(axireqArb_io_in_21_bits_entryid),
    .io_in_21_bits_arid(axireqArb_io_in_21_bits_arid),
    .io_in_21_bits_ardata(axireqArb_io_in_21_bits_ardata),
    .io_in_21_bits_respStatus(axireqArb_io_in_21_bits_respStatus),
    .io_in_21_bits_rsize(axireqArb_io_in_21_bits_rsize),
    .io_in_22_valid(axireqArb_io_in_22_valid),
    .io_in_22_bits_raddress(axireqArb_io_in_22_bits_raddress),
    .io_in_22_bits_entryid(axireqArb_io_in_22_bits_entryid),
    .io_in_22_bits_arid(axireqArb_io_in_22_bits_arid),
    .io_in_22_bits_ardata(axireqArb_io_in_22_bits_ardata),
    .io_in_22_bits_respStatus(axireqArb_io_in_22_bits_respStatus),
    .io_in_22_bits_rsize(axireqArb_io_in_22_bits_rsize),
    .io_in_23_valid(axireqArb_io_in_23_valid),
    .io_in_23_bits_raddress(axireqArb_io_in_23_bits_raddress),
    .io_in_23_bits_entryid(axireqArb_io_in_23_bits_entryid),
    .io_in_23_bits_arid(axireqArb_io_in_23_bits_arid),
    .io_in_23_bits_ardata(axireqArb_io_in_23_bits_ardata),
    .io_in_23_bits_respStatus(axireqArb_io_in_23_bits_respStatus),
    .io_in_23_bits_rsize(axireqArb_io_in_23_bits_rsize),
    .io_in_24_valid(axireqArb_io_in_24_valid),
    .io_in_24_bits_raddress(axireqArb_io_in_24_bits_raddress),
    .io_in_24_bits_entryid(axireqArb_io_in_24_bits_entryid),
    .io_in_24_bits_arid(axireqArb_io_in_24_bits_arid),
    .io_in_24_bits_ardata(axireqArb_io_in_24_bits_ardata),
    .io_in_24_bits_respStatus(axireqArb_io_in_24_bits_respStatus),
    .io_in_24_bits_rsize(axireqArb_io_in_24_bits_rsize),
    .io_in_25_valid(axireqArb_io_in_25_valid),
    .io_in_25_bits_raddress(axireqArb_io_in_25_bits_raddress),
    .io_in_25_bits_entryid(axireqArb_io_in_25_bits_entryid),
    .io_in_25_bits_arid(axireqArb_io_in_25_bits_arid),
    .io_in_25_bits_ardata(axireqArb_io_in_25_bits_ardata),
    .io_in_25_bits_respStatus(axireqArb_io_in_25_bits_respStatus),
    .io_in_25_bits_rsize(axireqArb_io_in_25_bits_rsize),
    .io_in_26_valid(axireqArb_io_in_26_valid),
    .io_in_26_bits_raddress(axireqArb_io_in_26_bits_raddress),
    .io_in_26_bits_entryid(axireqArb_io_in_26_bits_entryid),
    .io_in_26_bits_arid(axireqArb_io_in_26_bits_arid),
    .io_in_26_bits_ardata(axireqArb_io_in_26_bits_ardata),
    .io_in_26_bits_respStatus(axireqArb_io_in_26_bits_respStatus),
    .io_in_26_bits_rsize(axireqArb_io_in_26_bits_rsize),
    .io_in_27_valid(axireqArb_io_in_27_valid),
    .io_in_27_bits_raddress(axireqArb_io_in_27_bits_raddress),
    .io_in_27_bits_entryid(axireqArb_io_in_27_bits_entryid),
    .io_in_27_bits_arid(axireqArb_io_in_27_bits_arid),
    .io_in_27_bits_ardata(axireqArb_io_in_27_bits_ardata),
    .io_in_27_bits_respStatus(axireqArb_io_in_27_bits_respStatus),
    .io_in_27_bits_rsize(axireqArb_io_in_27_bits_rsize),
    .io_in_28_valid(axireqArb_io_in_28_valid),
    .io_in_28_bits_raddress(axireqArb_io_in_28_bits_raddress),
    .io_in_28_bits_entryid(axireqArb_io_in_28_bits_entryid),
    .io_in_28_bits_arid(axireqArb_io_in_28_bits_arid),
    .io_in_28_bits_ardata(axireqArb_io_in_28_bits_ardata),
    .io_in_28_bits_respStatus(axireqArb_io_in_28_bits_respStatus),
    .io_in_28_bits_rsize(axireqArb_io_in_28_bits_rsize),
    .io_in_29_valid(axireqArb_io_in_29_valid),
    .io_in_29_bits_raddress(axireqArb_io_in_29_bits_raddress),
    .io_in_29_bits_entryid(axireqArb_io_in_29_bits_entryid),
    .io_in_29_bits_arid(axireqArb_io_in_29_bits_arid),
    .io_in_29_bits_ardata(axireqArb_io_in_29_bits_ardata),
    .io_in_29_bits_respStatus(axireqArb_io_in_29_bits_respStatus),
    .io_in_29_bits_rsize(axireqArb_io_in_29_bits_rsize),
    .io_in_30_valid(axireqArb_io_in_30_valid),
    .io_in_30_bits_raddress(axireqArb_io_in_30_bits_raddress),
    .io_in_30_bits_entryid(axireqArb_io_in_30_bits_entryid),
    .io_in_30_bits_arid(axireqArb_io_in_30_bits_arid),
    .io_in_30_bits_ardata(axireqArb_io_in_30_bits_ardata),
    .io_in_30_bits_respStatus(axireqArb_io_in_30_bits_respStatus),
    .io_in_30_bits_rsize(axireqArb_io_in_30_bits_rsize),
    .io_in_31_valid(axireqArb_io_in_31_valid),
    .io_in_31_bits_raddress(axireqArb_io_in_31_bits_raddress),
    .io_in_31_bits_entryid(axireqArb_io_in_31_bits_entryid),
    .io_in_31_bits_arid(axireqArb_io_in_31_bits_arid),
    .io_in_31_bits_ardata(axireqArb_io_in_31_bits_ardata),
    .io_in_31_bits_respStatus(axireqArb_io_in_31_bits_respStatus),
    .io_in_31_bits_rsize(axireqArb_io_in_31_bits_rsize),
    .io_out_valid(axireqArb_io_out_valid),
    .io_out_bits_raddress(axireqArb_io_out_bits_raddress),
    .io_out_bits_entryid(axireqArb_io_out_bits_entryid),
    .io_out_bits_arid(axireqArb_io_out_bits_arid),
    .io_out_bits_ardata(axireqArb_io_out_bits_ardata),
    .io_out_bits_respStatus(axireqArb_io_out_bits_respStatus),
    .io_out_bits_rsize(axireqArb_io_out_bits_rsize),
    .io_chosen(axireqArb_io_chosen)
  );
  Arbiter axirespArb ( // @[ReadStack.scala 66:26]
    .io_in_0_valid(axirespArb_io_in_0_valid),
    .io_in_0_bits_raddress(axirespArb_io_in_0_bits_raddress),
    .io_in_0_bits_entryid(axirespArb_io_in_0_bits_entryid),
    .io_in_0_bits_arid(axirespArb_io_in_0_bits_arid),
    .io_in_0_bits_ardata(axirespArb_io_in_0_bits_ardata),
    .io_in_0_bits_respStatus(axirespArb_io_in_0_bits_respStatus),
    .io_in_0_bits_rsize(axirespArb_io_in_0_bits_rsize),
    .io_in_1_valid(axirespArb_io_in_1_valid),
    .io_in_1_bits_raddress(axirespArb_io_in_1_bits_raddress),
    .io_in_1_bits_entryid(axirespArb_io_in_1_bits_entryid),
    .io_in_1_bits_arid(axirespArb_io_in_1_bits_arid),
    .io_in_1_bits_ardata(axirespArb_io_in_1_bits_ardata),
    .io_in_1_bits_respStatus(axirespArb_io_in_1_bits_respStatus),
    .io_in_1_bits_rsize(axirespArb_io_in_1_bits_rsize),
    .io_in_2_valid(axirespArb_io_in_2_valid),
    .io_in_2_bits_raddress(axirespArb_io_in_2_bits_raddress),
    .io_in_2_bits_entryid(axirespArb_io_in_2_bits_entryid),
    .io_in_2_bits_arid(axirespArb_io_in_2_bits_arid),
    .io_in_2_bits_ardata(axirespArb_io_in_2_bits_ardata),
    .io_in_2_bits_respStatus(axirespArb_io_in_2_bits_respStatus),
    .io_in_2_bits_rsize(axirespArb_io_in_2_bits_rsize),
    .io_in_3_valid(axirespArb_io_in_3_valid),
    .io_in_3_bits_raddress(axirespArb_io_in_3_bits_raddress),
    .io_in_3_bits_entryid(axirespArb_io_in_3_bits_entryid),
    .io_in_3_bits_arid(axirespArb_io_in_3_bits_arid),
    .io_in_3_bits_ardata(axirespArb_io_in_3_bits_ardata),
    .io_in_3_bits_respStatus(axirespArb_io_in_3_bits_respStatus),
    .io_in_3_bits_rsize(axirespArb_io_in_3_bits_rsize),
    .io_in_4_valid(axirespArb_io_in_4_valid),
    .io_in_4_bits_raddress(axirespArb_io_in_4_bits_raddress),
    .io_in_4_bits_entryid(axirespArb_io_in_4_bits_entryid),
    .io_in_4_bits_arid(axirespArb_io_in_4_bits_arid),
    .io_in_4_bits_ardata(axirespArb_io_in_4_bits_ardata),
    .io_in_4_bits_respStatus(axirespArb_io_in_4_bits_respStatus),
    .io_in_4_bits_rsize(axirespArb_io_in_4_bits_rsize),
    .io_in_5_valid(axirespArb_io_in_5_valid),
    .io_in_5_bits_raddress(axirespArb_io_in_5_bits_raddress),
    .io_in_5_bits_entryid(axirespArb_io_in_5_bits_entryid),
    .io_in_5_bits_arid(axirespArb_io_in_5_bits_arid),
    .io_in_5_bits_ardata(axirespArb_io_in_5_bits_ardata),
    .io_in_5_bits_respStatus(axirespArb_io_in_5_bits_respStatus),
    .io_in_5_bits_rsize(axirespArb_io_in_5_bits_rsize),
    .io_in_6_valid(axirespArb_io_in_6_valid),
    .io_in_6_bits_raddress(axirespArb_io_in_6_bits_raddress),
    .io_in_6_bits_entryid(axirespArb_io_in_6_bits_entryid),
    .io_in_6_bits_arid(axirespArb_io_in_6_bits_arid),
    .io_in_6_bits_ardata(axirespArb_io_in_6_bits_ardata),
    .io_in_6_bits_respStatus(axirespArb_io_in_6_bits_respStatus),
    .io_in_6_bits_rsize(axirespArb_io_in_6_bits_rsize),
    .io_in_7_valid(axirespArb_io_in_7_valid),
    .io_in_7_bits_raddress(axirespArb_io_in_7_bits_raddress),
    .io_in_7_bits_entryid(axirespArb_io_in_7_bits_entryid),
    .io_in_7_bits_arid(axirespArb_io_in_7_bits_arid),
    .io_in_7_bits_ardata(axirespArb_io_in_7_bits_ardata),
    .io_in_7_bits_respStatus(axirespArb_io_in_7_bits_respStatus),
    .io_in_7_bits_rsize(axirespArb_io_in_7_bits_rsize),
    .io_in_8_valid(axirespArb_io_in_8_valid),
    .io_in_8_bits_raddress(axirespArb_io_in_8_bits_raddress),
    .io_in_8_bits_entryid(axirespArb_io_in_8_bits_entryid),
    .io_in_8_bits_arid(axirespArb_io_in_8_bits_arid),
    .io_in_8_bits_ardata(axirespArb_io_in_8_bits_ardata),
    .io_in_8_bits_respStatus(axirespArb_io_in_8_bits_respStatus),
    .io_in_8_bits_rsize(axirespArb_io_in_8_bits_rsize),
    .io_in_9_valid(axirespArb_io_in_9_valid),
    .io_in_9_bits_raddress(axirespArb_io_in_9_bits_raddress),
    .io_in_9_bits_entryid(axirespArb_io_in_9_bits_entryid),
    .io_in_9_bits_arid(axirespArb_io_in_9_bits_arid),
    .io_in_9_bits_ardata(axirespArb_io_in_9_bits_ardata),
    .io_in_9_bits_respStatus(axirespArb_io_in_9_bits_respStatus),
    .io_in_9_bits_rsize(axirespArb_io_in_9_bits_rsize),
    .io_in_10_valid(axirespArb_io_in_10_valid),
    .io_in_10_bits_raddress(axirespArb_io_in_10_bits_raddress),
    .io_in_10_bits_entryid(axirespArb_io_in_10_bits_entryid),
    .io_in_10_bits_arid(axirespArb_io_in_10_bits_arid),
    .io_in_10_bits_ardata(axirespArb_io_in_10_bits_ardata),
    .io_in_10_bits_respStatus(axirespArb_io_in_10_bits_respStatus),
    .io_in_10_bits_rsize(axirespArb_io_in_10_bits_rsize),
    .io_in_11_valid(axirespArb_io_in_11_valid),
    .io_in_11_bits_raddress(axirespArb_io_in_11_bits_raddress),
    .io_in_11_bits_entryid(axirespArb_io_in_11_bits_entryid),
    .io_in_11_bits_arid(axirespArb_io_in_11_bits_arid),
    .io_in_11_bits_ardata(axirespArb_io_in_11_bits_ardata),
    .io_in_11_bits_respStatus(axirespArb_io_in_11_bits_respStatus),
    .io_in_11_bits_rsize(axirespArb_io_in_11_bits_rsize),
    .io_in_12_valid(axirespArb_io_in_12_valid),
    .io_in_12_bits_raddress(axirespArb_io_in_12_bits_raddress),
    .io_in_12_bits_entryid(axirespArb_io_in_12_bits_entryid),
    .io_in_12_bits_arid(axirespArb_io_in_12_bits_arid),
    .io_in_12_bits_ardata(axirespArb_io_in_12_bits_ardata),
    .io_in_12_bits_respStatus(axirespArb_io_in_12_bits_respStatus),
    .io_in_12_bits_rsize(axirespArb_io_in_12_bits_rsize),
    .io_in_13_valid(axirespArb_io_in_13_valid),
    .io_in_13_bits_raddress(axirespArb_io_in_13_bits_raddress),
    .io_in_13_bits_entryid(axirespArb_io_in_13_bits_entryid),
    .io_in_13_bits_arid(axirespArb_io_in_13_bits_arid),
    .io_in_13_bits_ardata(axirespArb_io_in_13_bits_ardata),
    .io_in_13_bits_respStatus(axirespArb_io_in_13_bits_respStatus),
    .io_in_13_bits_rsize(axirespArb_io_in_13_bits_rsize),
    .io_in_14_valid(axirespArb_io_in_14_valid),
    .io_in_14_bits_raddress(axirespArb_io_in_14_bits_raddress),
    .io_in_14_bits_entryid(axirespArb_io_in_14_bits_entryid),
    .io_in_14_bits_arid(axirespArb_io_in_14_bits_arid),
    .io_in_14_bits_ardata(axirespArb_io_in_14_bits_ardata),
    .io_in_14_bits_respStatus(axirespArb_io_in_14_bits_respStatus),
    .io_in_14_bits_rsize(axirespArb_io_in_14_bits_rsize),
    .io_in_15_valid(axirespArb_io_in_15_valid),
    .io_in_15_bits_raddress(axirespArb_io_in_15_bits_raddress),
    .io_in_15_bits_entryid(axirespArb_io_in_15_bits_entryid),
    .io_in_15_bits_arid(axirespArb_io_in_15_bits_arid),
    .io_in_15_bits_ardata(axirespArb_io_in_15_bits_ardata),
    .io_in_15_bits_respStatus(axirespArb_io_in_15_bits_respStatus),
    .io_in_15_bits_rsize(axirespArb_io_in_15_bits_rsize),
    .io_in_16_valid(axirespArb_io_in_16_valid),
    .io_in_16_bits_raddress(axirespArb_io_in_16_bits_raddress),
    .io_in_16_bits_entryid(axirespArb_io_in_16_bits_entryid),
    .io_in_16_bits_arid(axirespArb_io_in_16_bits_arid),
    .io_in_16_bits_ardata(axirespArb_io_in_16_bits_ardata),
    .io_in_16_bits_respStatus(axirespArb_io_in_16_bits_respStatus),
    .io_in_16_bits_rsize(axirespArb_io_in_16_bits_rsize),
    .io_in_17_valid(axirespArb_io_in_17_valid),
    .io_in_17_bits_raddress(axirespArb_io_in_17_bits_raddress),
    .io_in_17_bits_entryid(axirespArb_io_in_17_bits_entryid),
    .io_in_17_bits_arid(axirespArb_io_in_17_bits_arid),
    .io_in_17_bits_ardata(axirespArb_io_in_17_bits_ardata),
    .io_in_17_bits_respStatus(axirespArb_io_in_17_bits_respStatus),
    .io_in_17_bits_rsize(axirespArb_io_in_17_bits_rsize),
    .io_in_18_valid(axirespArb_io_in_18_valid),
    .io_in_18_bits_raddress(axirespArb_io_in_18_bits_raddress),
    .io_in_18_bits_entryid(axirespArb_io_in_18_bits_entryid),
    .io_in_18_bits_arid(axirespArb_io_in_18_bits_arid),
    .io_in_18_bits_ardata(axirespArb_io_in_18_bits_ardata),
    .io_in_18_bits_respStatus(axirespArb_io_in_18_bits_respStatus),
    .io_in_18_bits_rsize(axirespArb_io_in_18_bits_rsize),
    .io_in_19_valid(axirespArb_io_in_19_valid),
    .io_in_19_bits_raddress(axirespArb_io_in_19_bits_raddress),
    .io_in_19_bits_entryid(axirespArb_io_in_19_bits_entryid),
    .io_in_19_bits_arid(axirespArb_io_in_19_bits_arid),
    .io_in_19_bits_ardata(axirespArb_io_in_19_bits_ardata),
    .io_in_19_bits_respStatus(axirespArb_io_in_19_bits_respStatus),
    .io_in_19_bits_rsize(axirespArb_io_in_19_bits_rsize),
    .io_in_20_valid(axirespArb_io_in_20_valid),
    .io_in_20_bits_raddress(axirespArb_io_in_20_bits_raddress),
    .io_in_20_bits_entryid(axirespArb_io_in_20_bits_entryid),
    .io_in_20_bits_arid(axirespArb_io_in_20_bits_arid),
    .io_in_20_bits_ardata(axirespArb_io_in_20_bits_ardata),
    .io_in_20_bits_respStatus(axirespArb_io_in_20_bits_respStatus),
    .io_in_20_bits_rsize(axirespArb_io_in_20_bits_rsize),
    .io_in_21_valid(axirespArb_io_in_21_valid),
    .io_in_21_bits_raddress(axirespArb_io_in_21_bits_raddress),
    .io_in_21_bits_entryid(axirespArb_io_in_21_bits_entryid),
    .io_in_21_bits_arid(axirespArb_io_in_21_bits_arid),
    .io_in_21_bits_ardata(axirespArb_io_in_21_bits_ardata),
    .io_in_21_bits_respStatus(axirespArb_io_in_21_bits_respStatus),
    .io_in_21_bits_rsize(axirespArb_io_in_21_bits_rsize),
    .io_in_22_valid(axirespArb_io_in_22_valid),
    .io_in_22_bits_raddress(axirespArb_io_in_22_bits_raddress),
    .io_in_22_bits_entryid(axirespArb_io_in_22_bits_entryid),
    .io_in_22_bits_arid(axirespArb_io_in_22_bits_arid),
    .io_in_22_bits_ardata(axirespArb_io_in_22_bits_ardata),
    .io_in_22_bits_respStatus(axirespArb_io_in_22_bits_respStatus),
    .io_in_22_bits_rsize(axirespArb_io_in_22_bits_rsize),
    .io_in_23_valid(axirespArb_io_in_23_valid),
    .io_in_23_bits_raddress(axirespArb_io_in_23_bits_raddress),
    .io_in_23_bits_entryid(axirespArb_io_in_23_bits_entryid),
    .io_in_23_bits_arid(axirespArb_io_in_23_bits_arid),
    .io_in_23_bits_ardata(axirespArb_io_in_23_bits_ardata),
    .io_in_23_bits_respStatus(axirespArb_io_in_23_bits_respStatus),
    .io_in_23_bits_rsize(axirespArb_io_in_23_bits_rsize),
    .io_in_24_valid(axirespArb_io_in_24_valid),
    .io_in_24_bits_raddress(axirespArb_io_in_24_bits_raddress),
    .io_in_24_bits_entryid(axirespArb_io_in_24_bits_entryid),
    .io_in_24_bits_arid(axirespArb_io_in_24_bits_arid),
    .io_in_24_bits_ardata(axirespArb_io_in_24_bits_ardata),
    .io_in_24_bits_respStatus(axirespArb_io_in_24_bits_respStatus),
    .io_in_24_bits_rsize(axirespArb_io_in_24_bits_rsize),
    .io_in_25_valid(axirespArb_io_in_25_valid),
    .io_in_25_bits_raddress(axirespArb_io_in_25_bits_raddress),
    .io_in_25_bits_entryid(axirespArb_io_in_25_bits_entryid),
    .io_in_25_bits_arid(axirespArb_io_in_25_bits_arid),
    .io_in_25_bits_ardata(axirespArb_io_in_25_bits_ardata),
    .io_in_25_bits_respStatus(axirespArb_io_in_25_bits_respStatus),
    .io_in_25_bits_rsize(axirespArb_io_in_25_bits_rsize),
    .io_in_26_valid(axirespArb_io_in_26_valid),
    .io_in_26_bits_raddress(axirespArb_io_in_26_bits_raddress),
    .io_in_26_bits_entryid(axirespArb_io_in_26_bits_entryid),
    .io_in_26_bits_arid(axirespArb_io_in_26_bits_arid),
    .io_in_26_bits_ardata(axirespArb_io_in_26_bits_ardata),
    .io_in_26_bits_respStatus(axirespArb_io_in_26_bits_respStatus),
    .io_in_26_bits_rsize(axirespArb_io_in_26_bits_rsize),
    .io_in_27_valid(axirespArb_io_in_27_valid),
    .io_in_27_bits_raddress(axirespArb_io_in_27_bits_raddress),
    .io_in_27_bits_entryid(axirespArb_io_in_27_bits_entryid),
    .io_in_27_bits_arid(axirespArb_io_in_27_bits_arid),
    .io_in_27_bits_ardata(axirespArb_io_in_27_bits_ardata),
    .io_in_27_bits_respStatus(axirespArb_io_in_27_bits_respStatus),
    .io_in_27_bits_rsize(axirespArb_io_in_27_bits_rsize),
    .io_in_28_valid(axirespArb_io_in_28_valid),
    .io_in_28_bits_raddress(axirespArb_io_in_28_bits_raddress),
    .io_in_28_bits_entryid(axirespArb_io_in_28_bits_entryid),
    .io_in_28_bits_arid(axirespArb_io_in_28_bits_arid),
    .io_in_28_bits_ardata(axirespArb_io_in_28_bits_ardata),
    .io_in_28_bits_respStatus(axirespArb_io_in_28_bits_respStatus),
    .io_in_28_bits_rsize(axirespArb_io_in_28_bits_rsize),
    .io_in_29_valid(axirespArb_io_in_29_valid),
    .io_in_29_bits_raddress(axirespArb_io_in_29_bits_raddress),
    .io_in_29_bits_entryid(axirespArb_io_in_29_bits_entryid),
    .io_in_29_bits_arid(axirespArb_io_in_29_bits_arid),
    .io_in_29_bits_ardata(axirespArb_io_in_29_bits_ardata),
    .io_in_29_bits_respStatus(axirespArb_io_in_29_bits_respStatus),
    .io_in_29_bits_rsize(axirespArb_io_in_29_bits_rsize),
    .io_in_30_valid(axirespArb_io_in_30_valid),
    .io_in_30_bits_raddress(axirespArb_io_in_30_bits_raddress),
    .io_in_30_bits_entryid(axirespArb_io_in_30_bits_entryid),
    .io_in_30_bits_arid(axirespArb_io_in_30_bits_arid),
    .io_in_30_bits_ardata(axirespArb_io_in_30_bits_ardata),
    .io_in_30_bits_respStatus(axirespArb_io_in_30_bits_respStatus),
    .io_in_30_bits_rsize(axirespArb_io_in_30_bits_rsize),
    .io_in_31_valid(axirespArb_io_in_31_valid),
    .io_in_31_bits_raddress(axirespArb_io_in_31_bits_raddress),
    .io_in_31_bits_entryid(axirespArb_io_in_31_bits_entryid),
    .io_in_31_bits_arid(axirespArb_io_in_31_bits_arid),
    .io_in_31_bits_ardata(axirespArb_io_in_31_bits_ardata),
    .io_in_31_bits_respStatus(axirespArb_io_in_31_bits_respStatus),
    .io_in_31_bits_rsize(axirespArb_io_in_31_bits_rsize),
    .io_out_valid(axirespArb_io_out_valid),
    .io_out_bits_raddress(axirespArb_io_out_bits_raddress),
    .io_out_bits_entryid(axirespArb_io_out_bits_entryid),
    .io_out_bits_arid(axirespArb_io_out_bits_arid),
    .io_out_bits_ardata(axirespArb_io_out_bits_ardata),
    .io_out_bits_respStatus(axirespArb_io_out_bits_respStatus),
    .io_out_bits_rsize(axirespArb_io_out_bits_rsize),
    .io_chosen(axirespArb_io_chosen)
  );
  assign io_axiReq_in_ar_ready = ~full; // @[ReadStack.scala 73:28]
  assign io_tlResp_in_d_ready = |_canReceive_T_64; // @[ReadStack.scala 150:82]
  assign io_tlReq_out_a_valid = axireqArb_io_out_valid; // @[ReadStack.scala 108:24]
  assign io_tlReq_out_a_bits_opcode = 3'h4; // @[ReadStack.scala 109:30]
  assign io_tlReq_out_a_bits_param = 3'h0; // @[ReadStack.scala 110:29]
  assign io_tlReq_out_a_bits_size = axireqArb_io_out_bits_rsize[2:0]; // @[ReadStack.scala 111:28]
  assign io_tlReq_out_a_bits_source = {axireqArb_io_out_bits_entryid,axireqArb_io_out_bits_arid}; // @[Cat.scala 31:58]
  assign io_tlReq_out_a_bits_address = axireqArb_io_out_bits_raddress; // @[ReadStack.scala 113:31]
  assign io_tlReq_out_a_bits_mask = {{24'd0}, _io_tlReq_out_a_bits_mask_T_1}; // @[ReadStack.scala 114:28]
  assign io_tlReq_out_a_bits_data = 256'h0; // @[ReadStack.scala 115:28]
  assign io_tlReq_out_a_bits_corrupt = 1'h0; // @[ReadStack.scala 116:31]
  assign io_axiResp_out_r_valid = axirespArb_io_out_valid; // @[ReadStack.scala 167:26]
  assign io_axiResp_out_r_bits_id = axirespArb_io_out_bits_arid; // @[ReadStack.scala 169:28]
  assign io_axiResp_out_r_bits_data = axirespArb_io_out_bits_ardata; // @[ReadStack.scala 168:30]
  assign io_axiResp_out_r_bits_resp = axirespArb_io_out_bits_respStatus[1:0]; // @[ReadStack.scala 170:30]
  assign io_axiResp_out_r_bits_last = 1'h1; // @[ReadStack.scala 174:30]
  assign axireqArb_io_in_0_valid = readStack_0_rvalid & _hasWaitTLReq_T & readStack_0_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_0_bits_raddress = readStack_0_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_0_bits_entryid = readStack_0_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_0_bits_arid = readStack_0_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_0_bits_ardata = readStack_0_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_0_bits_respStatus = readStack_0_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_0_bits_rsize = readStack_0_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_valid = readStack_1_rvalid & _hasWaitTLReq_T_1 & readStack_1_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_1_bits_raddress = readStack_1_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_bits_entryid = readStack_1_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_bits_arid = readStack_1_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_bits_ardata = readStack_1_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_bits_respStatus = readStack_1_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_1_bits_rsize = readStack_1_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_valid = readStack_2_rvalid & _hasWaitTLReq_T_2 & readStack_2_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_2_bits_raddress = readStack_2_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_bits_entryid = readStack_2_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_bits_arid = readStack_2_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_bits_ardata = readStack_2_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_bits_respStatus = readStack_2_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_2_bits_rsize = readStack_2_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_valid = readStack_3_rvalid & _hasWaitTLReq_T_3 & readStack_3_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_3_bits_raddress = readStack_3_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_bits_entryid = readStack_3_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_bits_arid = readStack_3_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_bits_ardata = readStack_3_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_bits_respStatus = readStack_3_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_3_bits_rsize = readStack_3_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_valid = readStack_4_rvalid & _hasWaitTLReq_T_4 & readStack_4_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_4_bits_raddress = readStack_4_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_bits_entryid = readStack_4_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_bits_arid = readStack_4_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_bits_ardata = readStack_4_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_bits_respStatus = readStack_4_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_4_bits_rsize = readStack_4_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_valid = readStack_5_rvalid & _hasWaitTLReq_T_5 & readStack_5_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_5_bits_raddress = readStack_5_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_bits_entryid = readStack_5_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_bits_arid = readStack_5_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_bits_ardata = readStack_5_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_bits_respStatus = readStack_5_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_5_bits_rsize = readStack_5_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_valid = readStack_6_rvalid & _hasWaitTLReq_T_6 & readStack_6_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_6_bits_raddress = readStack_6_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_bits_entryid = readStack_6_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_bits_arid = readStack_6_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_bits_ardata = readStack_6_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_bits_respStatus = readStack_6_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_6_bits_rsize = readStack_6_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_valid = readStack_7_rvalid & _hasWaitTLReq_T_7 & readStack_7_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_7_bits_raddress = readStack_7_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_bits_entryid = readStack_7_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_bits_arid = readStack_7_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_bits_ardata = readStack_7_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_bits_respStatus = readStack_7_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_7_bits_rsize = readStack_7_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_valid = readStack_8_rvalid & _hasWaitTLReq_T_8 & readStack_8_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_8_bits_raddress = readStack_8_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_bits_entryid = readStack_8_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_bits_arid = readStack_8_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_bits_ardata = readStack_8_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_bits_respStatus = readStack_8_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_8_bits_rsize = readStack_8_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_valid = readStack_9_rvalid & _hasWaitTLReq_T_9 & readStack_9_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_9_bits_raddress = readStack_9_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_bits_entryid = readStack_9_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_bits_arid = readStack_9_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_bits_ardata = readStack_9_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_bits_respStatus = readStack_9_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_9_bits_rsize = readStack_9_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_valid = readStack_10_rvalid & _hasWaitTLReq_T_10 & readStack_10_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_10_bits_raddress = readStack_10_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_bits_entryid = readStack_10_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_bits_arid = readStack_10_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_bits_ardata = readStack_10_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_bits_respStatus = readStack_10_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_10_bits_rsize = readStack_10_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_valid = readStack_11_rvalid & _hasWaitTLReq_T_11 & readStack_11_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_11_bits_raddress = readStack_11_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_bits_entryid = readStack_11_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_bits_arid = readStack_11_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_bits_ardata = readStack_11_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_bits_respStatus = readStack_11_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_11_bits_rsize = readStack_11_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_valid = readStack_12_rvalid & _hasWaitTLReq_T_12 & readStack_12_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_12_bits_raddress = readStack_12_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_bits_entryid = readStack_12_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_bits_arid = readStack_12_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_bits_ardata = readStack_12_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_bits_respStatus = readStack_12_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_12_bits_rsize = readStack_12_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_valid = readStack_13_rvalid & _hasWaitTLReq_T_13 & readStack_13_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_13_bits_raddress = readStack_13_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_bits_entryid = readStack_13_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_bits_arid = readStack_13_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_bits_ardata = readStack_13_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_bits_respStatus = readStack_13_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_13_bits_rsize = readStack_13_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_valid = readStack_14_rvalid & _hasWaitTLReq_T_14 & readStack_14_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_14_bits_raddress = readStack_14_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_bits_entryid = readStack_14_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_bits_arid = readStack_14_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_bits_ardata = readStack_14_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_bits_respStatus = readStack_14_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_14_bits_rsize = readStack_14_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_valid = readStack_15_rvalid & _hasWaitTLReq_T_15 & readStack_15_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_15_bits_raddress = readStack_15_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_bits_entryid = readStack_15_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_bits_arid = readStack_15_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_bits_ardata = readStack_15_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_bits_respStatus = readStack_15_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_15_bits_rsize = readStack_15_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_valid = readStack_16_rvalid & _hasWaitTLReq_T_16 & readStack_16_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_16_bits_raddress = readStack_16_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_bits_entryid = readStack_16_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_bits_arid = readStack_16_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_bits_ardata = readStack_16_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_bits_respStatus = readStack_16_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_16_bits_rsize = readStack_16_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_valid = readStack_17_rvalid & _hasWaitTLReq_T_17 & readStack_17_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_17_bits_raddress = readStack_17_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_bits_entryid = readStack_17_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_bits_arid = readStack_17_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_bits_ardata = readStack_17_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_bits_respStatus = readStack_17_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_17_bits_rsize = readStack_17_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_valid = readStack_18_rvalid & _hasWaitTLReq_T_18 & readStack_18_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_18_bits_raddress = readStack_18_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_bits_entryid = readStack_18_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_bits_arid = readStack_18_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_bits_ardata = readStack_18_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_bits_respStatus = readStack_18_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_18_bits_rsize = readStack_18_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_valid = readStack_19_rvalid & _hasWaitTLReq_T_19 & readStack_19_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_19_bits_raddress = readStack_19_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_bits_entryid = readStack_19_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_bits_arid = readStack_19_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_bits_ardata = readStack_19_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_bits_respStatus = readStack_19_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_19_bits_rsize = readStack_19_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_valid = readStack_20_rvalid & _hasWaitTLReq_T_20 & readStack_20_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_20_bits_raddress = readStack_20_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_bits_entryid = readStack_20_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_bits_arid = readStack_20_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_bits_ardata = readStack_20_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_bits_respStatus = readStack_20_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_20_bits_rsize = readStack_20_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_valid = readStack_21_rvalid & _hasWaitTLReq_T_21 & readStack_21_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_21_bits_raddress = readStack_21_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_bits_entryid = readStack_21_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_bits_arid = readStack_21_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_bits_ardata = readStack_21_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_bits_respStatus = readStack_21_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_21_bits_rsize = readStack_21_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_valid = readStack_22_rvalid & _hasWaitTLReq_T_22 & readStack_22_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_22_bits_raddress = readStack_22_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_bits_entryid = readStack_22_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_bits_arid = readStack_22_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_bits_ardata = readStack_22_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_bits_respStatus = readStack_22_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_22_bits_rsize = readStack_22_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_valid = readStack_23_rvalid & _hasWaitTLReq_T_23 & readStack_23_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_23_bits_raddress = readStack_23_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_bits_entryid = readStack_23_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_bits_arid = readStack_23_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_bits_ardata = readStack_23_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_bits_respStatus = readStack_23_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_23_bits_rsize = readStack_23_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_valid = readStack_24_rvalid & _hasWaitTLReq_T_24 & readStack_24_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_24_bits_raddress = readStack_24_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_bits_entryid = readStack_24_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_bits_arid = readStack_24_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_bits_ardata = readStack_24_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_bits_respStatus = readStack_24_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_24_bits_rsize = readStack_24_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_valid = readStack_25_rvalid & _hasWaitTLReq_T_25 & readStack_25_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_25_bits_raddress = readStack_25_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_bits_entryid = readStack_25_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_bits_arid = readStack_25_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_bits_ardata = readStack_25_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_bits_respStatus = readStack_25_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_25_bits_rsize = readStack_25_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_valid = readStack_26_rvalid & _hasWaitTLReq_T_26 & readStack_26_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_26_bits_raddress = readStack_26_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_bits_entryid = readStack_26_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_bits_arid = readStack_26_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_bits_ardata = readStack_26_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_bits_respStatus = readStack_26_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_26_bits_rsize = readStack_26_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_valid = readStack_27_rvalid & _hasWaitTLReq_T_27 & readStack_27_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_27_bits_raddress = readStack_27_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_bits_entryid = readStack_27_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_bits_arid = readStack_27_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_bits_ardata = readStack_27_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_bits_respStatus = readStack_27_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_27_bits_rsize = readStack_27_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_valid = readStack_28_rvalid & _hasWaitTLReq_T_28 & readStack_28_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_28_bits_raddress = readStack_28_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_bits_entryid = readStack_28_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_bits_arid = readStack_28_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_bits_ardata = readStack_28_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_bits_respStatus = readStack_28_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_28_bits_rsize = readStack_28_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_valid = readStack_29_rvalid & _hasWaitTLReq_T_29 & readStack_29_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_29_bits_raddress = readStack_29_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_bits_entryid = readStack_29_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_bits_arid = readStack_29_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_bits_ardata = readStack_29_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_bits_respStatus = readStack_29_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_29_bits_rsize = readStack_29_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_valid = readStack_30_rvalid & _hasWaitTLReq_T_30 & readStack_30_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_30_bits_raddress = readStack_30_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_bits_entryid = readStack_30_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_bits_arid = readStack_30_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_bits_ardata = readStack_30_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_bits_respStatus = readStack_30_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_30_bits_rsize = readStack_30_rsize; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_valid = readStack_31_rvalid & _hasWaitTLReq_T_31 & readStack_31_entryFifoId == 6'h0; // @[ReadStack.scala 104:59]
  assign axireqArb_io_in_31_bits_raddress = readStack_31_raddress; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_bits_entryid = readStack_31_entryid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_bits_arid = readStack_31_arid; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_bits_ardata = readStack_31_ardata; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_bits_respStatus = readStack_31_respStatus; // @[ReadStack.scala 105:15]
  assign axireqArb_io_in_31_bits_rsize = readStack_31_rsize; // @[ReadStack.scala 105:15]
  assign axirespArb_io_in_0_valid = _GEN_1184 == 3'h3 & readStack_0_rvalid & readStack_0_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_0_bits_raddress = readStack_0_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_0_bits_entryid = readStack_0_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_0_bits_arid = readStack_0_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_0_bits_ardata = readStack_0_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_0_bits_respStatus = readStack_0_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_0_bits_rsize = readStack_0_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_valid = _GEN_1185 == 3'h3 & readStack_1_rvalid & readStack_1_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_1_bits_raddress = readStack_1_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_bits_entryid = readStack_1_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_bits_arid = readStack_1_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_bits_ardata = readStack_1_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_bits_respStatus = readStack_1_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_1_bits_rsize = readStack_1_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_valid = _GEN_1186 == 3'h3 & readStack_2_rvalid & readStack_2_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_2_bits_raddress = readStack_2_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_bits_entryid = readStack_2_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_bits_arid = readStack_2_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_bits_ardata = readStack_2_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_bits_respStatus = readStack_2_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_2_bits_rsize = readStack_2_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_valid = _GEN_1187 == 3'h3 & readStack_3_rvalid & readStack_3_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_3_bits_raddress = readStack_3_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_bits_entryid = readStack_3_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_bits_arid = readStack_3_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_bits_ardata = readStack_3_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_bits_respStatus = readStack_3_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_3_bits_rsize = readStack_3_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_valid = _GEN_1188 == 3'h3 & readStack_4_rvalid & readStack_4_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_4_bits_raddress = readStack_4_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_bits_entryid = readStack_4_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_bits_arid = readStack_4_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_bits_ardata = readStack_4_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_bits_respStatus = readStack_4_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_4_bits_rsize = readStack_4_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_valid = _GEN_1189 == 3'h3 & readStack_5_rvalid & readStack_5_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_5_bits_raddress = readStack_5_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_bits_entryid = readStack_5_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_bits_arid = readStack_5_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_bits_ardata = readStack_5_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_bits_respStatus = readStack_5_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_5_bits_rsize = readStack_5_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_valid = _GEN_1190 == 3'h3 & readStack_6_rvalid & readStack_6_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_6_bits_raddress = readStack_6_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_bits_entryid = readStack_6_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_bits_arid = readStack_6_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_bits_ardata = readStack_6_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_bits_respStatus = readStack_6_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_6_bits_rsize = readStack_6_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_valid = _GEN_1191 == 3'h3 & readStack_7_rvalid & readStack_7_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_7_bits_raddress = readStack_7_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_bits_entryid = readStack_7_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_bits_arid = readStack_7_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_bits_ardata = readStack_7_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_bits_respStatus = readStack_7_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_7_bits_rsize = readStack_7_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_valid = _GEN_1192 == 3'h3 & readStack_8_rvalid & readStack_8_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_8_bits_raddress = readStack_8_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_bits_entryid = readStack_8_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_bits_arid = readStack_8_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_bits_ardata = readStack_8_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_bits_respStatus = readStack_8_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_8_bits_rsize = readStack_8_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_valid = _GEN_1193 == 3'h3 & readStack_9_rvalid & readStack_9_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_9_bits_raddress = readStack_9_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_bits_entryid = readStack_9_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_bits_arid = readStack_9_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_bits_ardata = readStack_9_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_bits_respStatus = readStack_9_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_9_bits_rsize = readStack_9_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_valid = _GEN_1194 == 3'h3 & readStack_10_rvalid & readStack_10_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_10_bits_raddress = readStack_10_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_bits_entryid = readStack_10_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_bits_arid = readStack_10_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_bits_ardata = readStack_10_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_bits_respStatus = readStack_10_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_10_bits_rsize = readStack_10_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_valid = _GEN_1195 == 3'h3 & readStack_11_rvalid & readStack_11_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_11_bits_raddress = readStack_11_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_bits_entryid = readStack_11_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_bits_arid = readStack_11_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_bits_ardata = readStack_11_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_bits_respStatus = readStack_11_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_11_bits_rsize = readStack_11_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_valid = _GEN_1196 == 3'h3 & readStack_12_rvalid & readStack_12_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_12_bits_raddress = readStack_12_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_bits_entryid = readStack_12_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_bits_arid = readStack_12_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_bits_ardata = readStack_12_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_bits_respStatus = readStack_12_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_12_bits_rsize = readStack_12_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_valid = _GEN_1197 == 3'h3 & readStack_13_rvalid & readStack_13_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_13_bits_raddress = readStack_13_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_bits_entryid = readStack_13_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_bits_arid = readStack_13_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_bits_ardata = readStack_13_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_bits_respStatus = readStack_13_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_13_bits_rsize = readStack_13_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_valid = _GEN_1198 == 3'h3 & readStack_14_rvalid & readStack_14_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_14_bits_raddress = readStack_14_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_bits_entryid = readStack_14_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_bits_arid = readStack_14_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_bits_ardata = readStack_14_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_bits_respStatus = readStack_14_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_14_bits_rsize = readStack_14_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_valid = _GEN_1199 == 3'h3 & readStack_15_rvalid & readStack_15_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_15_bits_raddress = readStack_15_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_bits_entryid = readStack_15_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_bits_arid = readStack_15_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_bits_ardata = readStack_15_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_bits_respStatus = readStack_15_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_15_bits_rsize = readStack_15_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_valid = _GEN_1200 == 3'h3 & readStack_16_rvalid & readStack_16_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_16_bits_raddress = readStack_16_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_bits_entryid = readStack_16_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_bits_arid = readStack_16_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_bits_ardata = readStack_16_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_bits_respStatus = readStack_16_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_16_bits_rsize = readStack_16_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_valid = _GEN_1201 == 3'h3 & readStack_17_rvalid & readStack_17_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_17_bits_raddress = readStack_17_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_bits_entryid = readStack_17_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_bits_arid = readStack_17_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_bits_ardata = readStack_17_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_bits_respStatus = readStack_17_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_17_bits_rsize = readStack_17_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_valid = _GEN_1202 == 3'h3 & readStack_18_rvalid & readStack_18_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_18_bits_raddress = readStack_18_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_bits_entryid = readStack_18_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_bits_arid = readStack_18_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_bits_ardata = readStack_18_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_bits_respStatus = readStack_18_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_18_bits_rsize = readStack_18_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_valid = _GEN_1203 == 3'h3 & readStack_19_rvalid & readStack_19_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_19_bits_raddress = readStack_19_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_bits_entryid = readStack_19_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_bits_arid = readStack_19_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_bits_ardata = readStack_19_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_bits_respStatus = readStack_19_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_19_bits_rsize = readStack_19_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_valid = _GEN_1204 == 3'h3 & readStack_20_rvalid & readStack_20_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_20_bits_raddress = readStack_20_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_bits_entryid = readStack_20_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_bits_arid = readStack_20_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_bits_ardata = readStack_20_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_bits_respStatus = readStack_20_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_20_bits_rsize = readStack_20_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_valid = _GEN_1205 == 3'h3 & readStack_21_rvalid & readStack_21_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_21_bits_raddress = readStack_21_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_bits_entryid = readStack_21_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_bits_arid = readStack_21_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_bits_ardata = readStack_21_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_bits_respStatus = readStack_21_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_21_bits_rsize = readStack_21_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_valid = _GEN_1206 == 3'h3 & readStack_22_rvalid & readStack_22_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_22_bits_raddress = readStack_22_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_bits_entryid = readStack_22_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_bits_arid = readStack_22_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_bits_ardata = readStack_22_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_bits_respStatus = readStack_22_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_22_bits_rsize = readStack_22_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_valid = _GEN_1207 == 3'h3 & readStack_23_rvalid & readStack_23_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_23_bits_raddress = readStack_23_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_bits_entryid = readStack_23_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_bits_arid = readStack_23_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_bits_ardata = readStack_23_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_bits_respStatus = readStack_23_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_23_bits_rsize = readStack_23_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_valid = _GEN_1208 == 3'h3 & readStack_24_rvalid & readStack_24_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_24_bits_raddress = readStack_24_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_bits_entryid = readStack_24_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_bits_arid = readStack_24_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_bits_ardata = readStack_24_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_bits_respStatus = readStack_24_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_24_bits_rsize = readStack_24_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_valid = _GEN_1209 == 3'h3 & readStack_25_rvalid & readStack_25_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_25_bits_raddress = readStack_25_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_bits_entryid = readStack_25_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_bits_arid = readStack_25_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_bits_ardata = readStack_25_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_bits_respStatus = readStack_25_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_25_bits_rsize = readStack_25_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_valid = _GEN_1210 == 3'h3 & readStack_26_rvalid & readStack_26_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_26_bits_raddress = readStack_26_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_bits_entryid = readStack_26_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_bits_arid = readStack_26_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_bits_ardata = readStack_26_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_bits_respStatus = readStack_26_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_26_bits_rsize = readStack_26_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_valid = _GEN_1211 == 3'h3 & readStack_27_rvalid & readStack_27_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_27_bits_raddress = readStack_27_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_bits_entryid = readStack_27_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_bits_arid = readStack_27_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_bits_ardata = readStack_27_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_bits_respStatus = readStack_27_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_27_bits_rsize = readStack_27_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_valid = _GEN_1212 == 3'h3 & readStack_28_rvalid & readStack_28_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_28_bits_raddress = readStack_28_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_bits_entryid = readStack_28_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_bits_arid = readStack_28_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_bits_ardata = readStack_28_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_bits_respStatus = readStack_28_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_28_bits_rsize = readStack_28_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_valid = _GEN_1213 == 3'h3 & readStack_29_rvalid & readStack_29_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_29_bits_raddress = readStack_29_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_bits_entryid = readStack_29_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_bits_arid = readStack_29_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_bits_ardata = readStack_29_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_bits_respStatus = readStack_29_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_29_bits_rsize = readStack_29_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_valid = _GEN_1214 == 3'h3 & readStack_30_rvalid & readStack_30_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_30_bits_raddress = readStack_30_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_bits_entryid = readStack_30_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_bits_arid = readStack_30_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_bits_ardata = readStack_30_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_bits_respStatus = readStack_30_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_30_bits_rsize = readStack_30_rsize; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_valid = _GEN_1215 == 3'h3 & readStack_31_rvalid & readStack_31_BeatFifoId == 6'h0; // @[ReadStack.scala 163:62]
  assign axirespArb_io_in_31_bits_raddress = readStack_31_raddress; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_bits_entryid = readStack_31_entryid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_bits_arid = readStack_31_arid; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_bits_ardata = readStack_31_ardata; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_bits_respStatus = readStack_31_respStatus; // @[ReadStack.scala 164:15]
  assign axirespArb_io_in_31_bits_rsize = readStack_31_rsize; // @[ReadStack.scala 164:15]
  always @(posedge clock) begin
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h0 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_0_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_0_rvalid <= _GEN_192;
      end
    end else begin
      readStack_0_rvalid <= _GEN_192;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h0 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_0_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h0 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_0_entryid <= _idxInsert_T_62;
        end else begin
          readStack_0_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h0 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_0_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h0 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_0_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h0 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_0_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h0 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_0_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_0_readStatus <= _GEN_320;
      end
    end else begin
      readStack_0_readStatus <= _GEN_320;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h0 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_0_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h0 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_0_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T & readStack_0_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_0_entryFifoId <= _readStack_0_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_0_entryFifoId <= _GEN_480;
      end
    end else begin
      readStack_0_entryFifoId <= _GEN_480;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_0_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_0_rvalid & readStack_0_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_0_BeatFifoId <= _readStack_0_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_0_BeatFifoId <= _GEN_896;
      end
    end else begin
      readStack_0_BeatFifoId <= _GEN_896;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_1_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_1_rvalid <= _GEN_193;
      end
    end else begin
      readStack_1_rvalid <= _GEN_193;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_1_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_1_entryid <= _idxInsert_T_62;
        end else begin
          readStack_1_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_1_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_1_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_1_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_1_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_1_readStatus <= _GEN_321;
      end
    end else begin
      readStack_1_readStatus <= _GEN_321;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_1_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_1_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_1 & readStack_1_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_1_entryFifoId <= _readStack_1_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_1_entryFifoId <= _GEN_481;
      end
    end else begin
      readStack_1_entryFifoId <= _GEN_481;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_1_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_1_rvalid & readStack_1_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_1_BeatFifoId <= _readStack_1_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_1_BeatFifoId <= _GEN_897;
      end
    end else begin
      readStack_1_BeatFifoId <= _GEN_897;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h2 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_2_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_2_rvalid <= _GEN_194;
      end
    end else begin
      readStack_2_rvalid <= _GEN_194;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h2 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_2_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h2 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_2_entryid <= _idxInsert_T_62;
        end else begin
          readStack_2_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h2 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_2_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h2 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_2_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h2 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_2_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h2 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_2_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_2_readStatus <= _GEN_322;
      end
    end else begin
      readStack_2_readStatus <= _GEN_322;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h2 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_2_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h2 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_2_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_2 & readStack_2_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_2_entryFifoId <= _readStack_2_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_2_entryFifoId <= _GEN_482;
      end
    end else begin
      readStack_2_entryFifoId <= _GEN_482;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_2_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_2_rvalid & readStack_2_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_2_BeatFifoId <= _readStack_2_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_2_BeatFifoId <= _GEN_898;
      end
    end else begin
      readStack_2_BeatFifoId <= _GEN_898;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h3 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_3_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_3_rvalid <= _GEN_195;
      end
    end else begin
      readStack_3_rvalid <= _GEN_195;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h3 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_3_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h3 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_3_entryid <= _idxInsert_T_62;
        end else begin
          readStack_3_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h3 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_3_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h3 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_3_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h3 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_3_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h3 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_3_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_3_readStatus <= _GEN_323;
      end
    end else begin
      readStack_3_readStatus <= _GEN_323;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h3 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_3_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h3 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_3_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_3 & readStack_3_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_3_entryFifoId <= _readStack_3_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_3_entryFifoId <= _GEN_483;
      end
    end else begin
      readStack_3_entryFifoId <= _GEN_483;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_3_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_3_rvalid & readStack_3_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_3_BeatFifoId <= _readStack_3_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_3_BeatFifoId <= _GEN_899;
      end
    end else begin
      readStack_3_BeatFifoId <= _GEN_899;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h4 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_4_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_4_rvalid <= _GEN_196;
      end
    end else begin
      readStack_4_rvalid <= _GEN_196;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h4 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_4_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h4 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_4_entryid <= _idxInsert_T_62;
        end else begin
          readStack_4_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h4 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_4_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h4 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_4_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h4 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_4_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h4 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_4_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_4_readStatus <= _GEN_324;
      end
    end else begin
      readStack_4_readStatus <= _GEN_324;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h4 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_4_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h4 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_4_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_4 & readStack_4_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_4_entryFifoId <= _readStack_4_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_4_entryFifoId <= _GEN_484;
      end
    end else begin
      readStack_4_entryFifoId <= _GEN_484;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_4_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_4_rvalid & readStack_4_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_4_BeatFifoId <= _readStack_4_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_4_BeatFifoId <= _GEN_900;
      end
    end else begin
      readStack_4_BeatFifoId <= _GEN_900;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h5 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_5_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_5_rvalid <= _GEN_197;
      end
    end else begin
      readStack_5_rvalid <= _GEN_197;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h5 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_5_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h5 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_5_entryid <= _idxInsert_T_62;
        end else begin
          readStack_5_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h5 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_5_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h5 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_5_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h5 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_5_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h5 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_5_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_5_readStatus <= _GEN_325;
      end
    end else begin
      readStack_5_readStatus <= _GEN_325;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h5 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_5_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h5 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_5_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_5 & readStack_5_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_5_entryFifoId <= _readStack_5_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_5_entryFifoId <= _GEN_485;
      end
    end else begin
      readStack_5_entryFifoId <= _GEN_485;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_5_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_5_rvalid & readStack_5_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_5_BeatFifoId <= _readStack_5_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_5_BeatFifoId <= _GEN_901;
      end
    end else begin
      readStack_5_BeatFifoId <= _GEN_901;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h6 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_6_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_6_rvalid <= _GEN_198;
      end
    end else begin
      readStack_6_rvalid <= _GEN_198;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h6 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_6_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h6 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_6_entryid <= _idxInsert_T_62;
        end else begin
          readStack_6_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h6 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_6_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h6 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_6_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h6 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_6_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h6 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_6_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_6_readStatus <= _GEN_326;
      end
    end else begin
      readStack_6_readStatus <= _GEN_326;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h6 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_6_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h6 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_6_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_6 & readStack_6_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_6_entryFifoId <= _readStack_6_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_6_entryFifoId <= _GEN_486;
      end
    end else begin
      readStack_6_entryFifoId <= _GEN_486;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_6_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_6_rvalid & readStack_6_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_6_BeatFifoId <= _readStack_6_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_6_BeatFifoId <= _GEN_902;
      end
    end else begin
      readStack_6_BeatFifoId <= _GEN_902;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h7 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_7_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_7_rvalid <= _GEN_199;
      end
    end else begin
      readStack_7_rvalid <= _GEN_199;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h7 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_7_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h7 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_7_entryid <= _idxInsert_T_62;
        end else begin
          readStack_7_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h7 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_7_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h7 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_7_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h7 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_7_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h7 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_7_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_7_readStatus <= _GEN_327;
      end
    end else begin
      readStack_7_readStatus <= _GEN_327;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h7 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_7_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h7 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_7_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_7 & readStack_7_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_7_entryFifoId <= _readStack_7_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_7_entryFifoId <= _GEN_487;
      end
    end else begin
      readStack_7_entryFifoId <= _GEN_487;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_7_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_7_rvalid & readStack_7_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_7_BeatFifoId <= _readStack_7_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_7_BeatFifoId <= _GEN_903;
      end
    end else begin
      readStack_7_BeatFifoId <= _GEN_903;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h8 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_8_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_8_rvalid <= _GEN_200;
      end
    end else begin
      readStack_8_rvalid <= _GEN_200;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h8 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_8_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h8 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_8_entryid <= _idxInsert_T_62;
        end else begin
          readStack_8_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h8 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_8_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h8 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_8_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h8 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_8_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h8 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_8_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_8_readStatus <= _GEN_328;
      end
    end else begin
      readStack_8_readStatus <= _GEN_328;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h8 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_8_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h8 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_8_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_8 & readStack_8_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_8_entryFifoId <= _readStack_8_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_8_entryFifoId <= _GEN_488;
      end
    end else begin
      readStack_8_entryFifoId <= _GEN_488;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_8_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_8_rvalid & readStack_8_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_8_BeatFifoId <= _readStack_8_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_8_BeatFifoId <= _GEN_904;
      end
    end else begin
      readStack_8_BeatFifoId <= _GEN_904;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h9 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_9_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_9_rvalid <= _GEN_201;
      end
    end else begin
      readStack_9_rvalid <= _GEN_201;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h9 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_9_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h9 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_9_entryid <= _idxInsert_T_62;
        end else begin
          readStack_9_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h9 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_9_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h9 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_9_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h9 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_9_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h9 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_9_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_9_readStatus <= _GEN_329;
      end
    end else begin
      readStack_9_readStatus <= _GEN_329;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h9 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_9_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h9 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_9_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_9 & readStack_9_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_9_entryFifoId <= _readStack_9_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_9_entryFifoId <= _GEN_489;
      end
    end else begin
      readStack_9_entryFifoId <= _GEN_489;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_9_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_9_rvalid & readStack_9_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_9_BeatFifoId <= _readStack_9_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_9_BeatFifoId <= _GEN_905;
      end
    end else begin
      readStack_9_BeatFifoId <= _GEN_905;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'ha == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_10_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_10_rvalid <= _GEN_202;
      end
    end else begin
      readStack_10_rvalid <= _GEN_202;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'ha == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_10_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'ha == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_10_entryid <= _idxInsert_T_62;
        end else begin
          readStack_10_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'ha == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_10_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'ha == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_10_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'ha == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_10_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'ha == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_10_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_10_readStatus <= _GEN_330;
      end
    end else begin
      readStack_10_readStatus <= _GEN_330;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'ha == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_10_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'ha == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_10_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_10 & readStack_10_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_10_entryFifoId <= _readStack_10_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_10_entryFifoId <= _GEN_490;
      end
    end else begin
      readStack_10_entryFifoId <= _GEN_490;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_10_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_10_rvalid & readStack_10_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_10_BeatFifoId <= _readStack_10_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_10_BeatFifoId <= _GEN_906;
      end
    end else begin
      readStack_10_BeatFifoId <= _GEN_906;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'hb == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_11_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_11_rvalid <= _GEN_203;
      end
    end else begin
      readStack_11_rvalid <= _GEN_203;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hb == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_11_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hb == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_11_entryid <= _idxInsert_T_62;
        end else begin
          readStack_11_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hb == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_11_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'hb == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_11_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'hb == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_11_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'hb == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_11_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_11_readStatus <= _GEN_331;
      end
    end else begin
      readStack_11_readStatus <= _GEN_331;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'hb == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_11_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hb == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_11_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_11 & readStack_11_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_11_entryFifoId <= _readStack_11_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_11_entryFifoId <= _GEN_491;
      end
    end else begin
      readStack_11_entryFifoId <= _GEN_491;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_11_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_11_rvalid & readStack_11_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_11_BeatFifoId <= _readStack_11_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_11_BeatFifoId <= _GEN_907;
      end
    end else begin
      readStack_11_BeatFifoId <= _GEN_907;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'hc == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_12_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_12_rvalid <= _GEN_204;
      end
    end else begin
      readStack_12_rvalid <= _GEN_204;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hc == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_12_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hc == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_12_entryid <= _idxInsert_T_62;
        end else begin
          readStack_12_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hc == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_12_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'hc == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_12_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'hc == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_12_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'hc == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_12_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_12_readStatus <= _GEN_332;
      end
    end else begin
      readStack_12_readStatus <= _GEN_332;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'hc == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_12_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hc == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_12_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_12 & readStack_12_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_12_entryFifoId <= _readStack_12_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_12_entryFifoId <= _GEN_492;
      end
    end else begin
      readStack_12_entryFifoId <= _GEN_492;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_12_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_12_rvalid & readStack_12_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_12_BeatFifoId <= _readStack_12_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_12_BeatFifoId <= _GEN_908;
      end
    end else begin
      readStack_12_BeatFifoId <= _GEN_908;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'hd == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_13_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_13_rvalid <= _GEN_205;
      end
    end else begin
      readStack_13_rvalid <= _GEN_205;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hd == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_13_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hd == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_13_entryid <= _idxInsert_T_62;
        end else begin
          readStack_13_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hd == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_13_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'hd == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_13_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'hd == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_13_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'hd == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_13_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_13_readStatus <= _GEN_333;
      end
    end else begin
      readStack_13_readStatus <= _GEN_333;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'hd == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_13_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hd == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_13_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_13 & readStack_13_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_13_entryFifoId <= _readStack_13_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_13_entryFifoId <= _GEN_493;
      end
    end else begin
      readStack_13_entryFifoId <= _GEN_493;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_13_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_13_rvalid & readStack_13_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_13_BeatFifoId <= _readStack_13_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_13_BeatFifoId <= _GEN_909;
      end
    end else begin
      readStack_13_BeatFifoId <= _GEN_909;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'he == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_14_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_14_rvalid <= _GEN_206;
      end
    end else begin
      readStack_14_rvalid <= _GEN_206;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'he == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_14_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'he == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_14_entryid <= _idxInsert_T_62;
        end else begin
          readStack_14_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'he == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_14_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'he == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_14_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'he == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_14_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'he == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_14_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_14_readStatus <= _GEN_334;
      end
    end else begin
      readStack_14_readStatus <= _GEN_334;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'he == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_14_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'he == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_14_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_14 & readStack_14_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_14_entryFifoId <= _readStack_14_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_14_entryFifoId <= _GEN_494;
      end
    end else begin
      readStack_14_entryFifoId <= _GEN_494;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_14_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_14_rvalid & readStack_14_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_14_BeatFifoId <= _readStack_14_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_14_BeatFifoId <= _GEN_910;
      end
    end else begin
      readStack_14_BeatFifoId <= _GEN_910;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'hf == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_15_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_15_rvalid <= _GEN_207;
      end
    end else begin
      readStack_15_rvalid <= _GEN_207;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hf == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_15_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hf == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_15_entryid <= _idxInsert_T_62;
        end else begin
          readStack_15_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hf == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_15_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'hf == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_15_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'hf == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_15_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'hf == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_15_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_15_readStatus <= _GEN_335;
      end
    end else begin
      readStack_15_readStatus <= _GEN_335;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'hf == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_15_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'hf == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_15_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_15 & readStack_15_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_15_entryFifoId <= _readStack_15_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_15_entryFifoId <= _GEN_495;
      end
    end else begin
      readStack_15_entryFifoId <= _GEN_495;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_15_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_15_rvalid & readStack_15_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_15_BeatFifoId <= _readStack_15_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_15_BeatFifoId <= _GEN_911;
      end
    end else begin
      readStack_15_BeatFifoId <= _GEN_911;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h10 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_16_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_16_rvalid <= _GEN_208;
      end
    end else begin
      readStack_16_rvalid <= _GEN_208;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h10 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_16_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h10 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_16_entryid <= _idxInsert_T_62;
        end else begin
          readStack_16_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h10 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_16_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h10 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_16_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h10 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_16_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h10 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_16_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_16_readStatus <= _GEN_336;
      end
    end else begin
      readStack_16_readStatus <= _GEN_336;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h10 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_16_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h10 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_16_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_16 & readStack_16_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_16_entryFifoId <= _readStack_16_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_16_entryFifoId <= _GEN_496;
      end
    end else begin
      readStack_16_entryFifoId <= _GEN_496;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_16_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_16_rvalid & readStack_16_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_16_BeatFifoId <= _readStack_16_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_16_BeatFifoId <= _GEN_912;
      end
    end else begin
      readStack_16_BeatFifoId <= _GEN_912;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h11 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_17_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_17_rvalid <= _GEN_209;
      end
    end else begin
      readStack_17_rvalid <= _GEN_209;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h11 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_17_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h11 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_17_entryid <= _idxInsert_T_62;
        end else begin
          readStack_17_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h11 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_17_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h11 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_17_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h11 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_17_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h11 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_17_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_17_readStatus <= _GEN_337;
      end
    end else begin
      readStack_17_readStatus <= _GEN_337;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h11 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_17_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h11 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_17_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_17 & readStack_17_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_17_entryFifoId <= _readStack_17_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_17_entryFifoId <= _GEN_497;
      end
    end else begin
      readStack_17_entryFifoId <= _GEN_497;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_17_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_17_rvalid & readStack_17_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_17_BeatFifoId <= _readStack_17_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_17_BeatFifoId <= _GEN_913;
      end
    end else begin
      readStack_17_BeatFifoId <= _GEN_913;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h12 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_18_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_18_rvalid <= _GEN_210;
      end
    end else begin
      readStack_18_rvalid <= _GEN_210;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h12 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_18_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h12 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_18_entryid <= _idxInsert_T_62;
        end else begin
          readStack_18_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h12 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_18_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h12 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_18_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h12 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_18_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h12 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_18_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_18_readStatus <= _GEN_338;
      end
    end else begin
      readStack_18_readStatus <= _GEN_338;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h12 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_18_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h12 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_18_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_18 & readStack_18_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_18_entryFifoId <= _readStack_18_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_18_entryFifoId <= _GEN_498;
      end
    end else begin
      readStack_18_entryFifoId <= _GEN_498;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_18_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_18_rvalid & readStack_18_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_18_BeatFifoId <= _readStack_18_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_18_BeatFifoId <= _GEN_914;
      end
    end else begin
      readStack_18_BeatFifoId <= _GEN_914;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h13 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_19_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_19_rvalid <= _GEN_211;
      end
    end else begin
      readStack_19_rvalid <= _GEN_211;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h13 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_19_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h13 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_19_entryid <= _idxInsert_T_62;
        end else begin
          readStack_19_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h13 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_19_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h13 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_19_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h13 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_19_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h13 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_19_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_19_readStatus <= _GEN_339;
      end
    end else begin
      readStack_19_readStatus <= _GEN_339;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h13 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_19_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h13 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_19_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_19 & readStack_19_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_19_entryFifoId <= _readStack_19_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_19_entryFifoId <= _GEN_499;
      end
    end else begin
      readStack_19_entryFifoId <= _GEN_499;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_19_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_19_rvalid & readStack_19_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_19_BeatFifoId <= _readStack_19_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_19_BeatFifoId <= _GEN_915;
      end
    end else begin
      readStack_19_BeatFifoId <= _GEN_915;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h14 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_20_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_20_rvalid <= _GEN_212;
      end
    end else begin
      readStack_20_rvalid <= _GEN_212;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h14 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_20_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h14 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_20_entryid <= _idxInsert_T_62;
        end else begin
          readStack_20_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h14 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_20_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h14 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_20_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h14 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_20_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h14 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_20_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_20_readStatus <= _GEN_340;
      end
    end else begin
      readStack_20_readStatus <= _GEN_340;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h14 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_20_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h14 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_20_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_20 & readStack_20_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_20_entryFifoId <= _readStack_20_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_20_entryFifoId <= _GEN_500;
      end
    end else begin
      readStack_20_entryFifoId <= _GEN_500;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_20_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_20_rvalid & readStack_20_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_20_BeatFifoId <= _readStack_20_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_20_BeatFifoId <= _GEN_916;
      end
    end else begin
      readStack_20_BeatFifoId <= _GEN_916;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h15 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_21_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_21_rvalid <= _GEN_213;
      end
    end else begin
      readStack_21_rvalid <= _GEN_213;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h15 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_21_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h15 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_21_entryid <= _idxInsert_T_62;
        end else begin
          readStack_21_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h15 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_21_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h15 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_21_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h15 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_21_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h15 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_21_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_21_readStatus <= _GEN_341;
      end
    end else begin
      readStack_21_readStatus <= _GEN_341;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h15 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_21_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h15 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_21_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_21 & readStack_21_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_21_entryFifoId <= _readStack_21_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_21_entryFifoId <= _GEN_501;
      end
    end else begin
      readStack_21_entryFifoId <= _GEN_501;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_21_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_21_rvalid & readStack_21_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_21_BeatFifoId <= _readStack_21_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_21_BeatFifoId <= _GEN_917;
      end
    end else begin
      readStack_21_BeatFifoId <= _GEN_917;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h16 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_22_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_22_rvalid <= _GEN_214;
      end
    end else begin
      readStack_22_rvalid <= _GEN_214;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h16 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_22_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h16 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_22_entryid <= _idxInsert_T_62;
        end else begin
          readStack_22_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h16 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_22_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h16 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_22_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h16 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_22_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h16 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_22_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_22_readStatus <= _GEN_342;
      end
    end else begin
      readStack_22_readStatus <= _GEN_342;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h16 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_22_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h16 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_22_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_22 & readStack_22_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_22_entryFifoId <= _readStack_22_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_22_entryFifoId <= _GEN_502;
      end
    end else begin
      readStack_22_entryFifoId <= _GEN_502;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_22_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_22_rvalid & readStack_22_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_22_BeatFifoId <= _readStack_22_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_22_BeatFifoId <= _GEN_918;
      end
    end else begin
      readStack_22_BeatFifoId <= _GEN_918;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h17 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_23_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_23_rvalid <= _GEN_215;
      end
    end else begin
      readStack_23_rvalid <= _GEN_215;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h17 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_23_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h17 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_23_entryid <= _idxInsert_T_62;
        end else begin
          readStack_23_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h17 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_23_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h17 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_23_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h17 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_23_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h17 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_23_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_23_readStatus <= _GEN_343;
      end
    end else begin
      readStack_23_readStatus <= _GEN_343;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h17 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_23_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h17 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_23_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_23 & readStack_23_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_23_entryFifoId <= _readStack_23_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_23_entryFifoId <= _GEN_503;
      end
    end else begin
      readStack_23_entryFifoId <= _GEN_503;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_23_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_23_rvalid & readStack_23_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_23_BeatFifoId <= _readStack_23_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_23_BeatFifoId <= _GEN_919;
      end
    end else begin
      readStack_23_BeatFifoId <= _GEN_919;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h18 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_24_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_24_rvalid <= _GEN_216;
      end
    end else begin
      readStack_24_rvalid <= _GEN_216;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h18 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_24_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h18 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_24_entryid <= _idxInsert_T_62;
        end else begin
          readStack_24_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h18 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_24_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h18 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_24_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h18 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_24_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h18 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_24_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_24_readStatus <= _GEN_344;
      end
    end else begin
      readStack_24_readStatus <= _GEN_344;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h18 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_24_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h18 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_24_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_24 & readStack_24_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_24_entryFifoId <= _readStack_24_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_24_entryFifoId <= _GEN_504;
      end
    end else begin
      readStack_24_entryFifoId <= _GEN_504;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_24_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_24_rvalid & readStack_24_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_24_BeatFifoId <= _readStack_24_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_24_BeatFifoId <= _GEN_920;
      end
    end else begin
      readStack_24_BeatFifoId <= _GEN_920;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h19 == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_25_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_25_rvalid <= _GEN_217;
      end
    end else begin
      readStack_25_rvalid <= _GEN_217;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h19 == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_25_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h19 == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_25_entryid <= _idxInsert_T_62;
        end else begin
          readStack_25_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h19 == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_25_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h19 == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_25_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h19 == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_25_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h19 == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_25_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_25_readStatus <= _GEN_345;
      end
    end else begin
      readStack_25_readStatus <= _GEN_345;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h19 == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_25_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h19 == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_25_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_25 & readStack_25_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_25_entryFifoId <= _readStack_25_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_25_entryFifoId <= _GEN_505;
      end
    end else begin
      readStack_25_entryFifoId <= _GEN_505;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_25_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_25_rvalid & readStack_25_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_25_BeatFifoId <= _readStack_25_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_25_BeatFifoId <= _GEN_921;
      end
    end else begin
      readStack_25_BeatFifoId <= _GEN_921;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1a == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_26_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_26_rvalid <= _GEN_218;
      end
    end else begin
      readStack_26_rvalid <= _GEN_218;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1a == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_26_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1a == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_26_entryid <= _idxInsert_T_62;
        end else begin
          readStack_26_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1a == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_26_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1a == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_26_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1a == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_26_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1a == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_26_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_26_readStatus <= _GEN_346;
      end
    end else begin
      readStack_26_readStatus <= _GEN_346;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1a == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_26_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1a == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_26_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_26 & readStack_26_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_26_entryFifoId <= _readStack_26_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_26_entryFifoId <= _GEN_506;
      end
    end else begin
      readStack_26_entryFifoId <= _GEN_506;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_26_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_26_rvalid & readStack_26_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_26_BeatFifoId <= _readStack_26_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_26_BeatFifoId <= _GEN_922;
      end
    end else begin
      readStack_26_BeatFifoId <= _GEN_922;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1b == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_27_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_27_rvalid <= _GEN_219;
      end
    end else begin
      readStack_27_rvalid <= _GEN_219;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1b == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_27_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1b == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_27_entryid <= _idxInsert_T_62;
        end else begin
          readStack_27_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1b == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_27_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1b == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_27_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1b == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_27_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1b == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_27_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_27_readStatus <= _GEN_347;
      end
    end else begin
      readStack_27_readStatus <= _GEN_347;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1b == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_27_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1b == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_27_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_27 & readStack_27_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_27_entryFifoId <= _readStack_27_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_27_entryFifoId <= _GEN_507;
      end
    end else begin
      readStack_27_entryFifoId <= _GEN_507;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_27_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_27_rvalid & readStack_27_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_27_BeatFifoId <= _readStack_27_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_27_BeatFifoId <= _GEN_923;
      end
    end else begin
      readStack_27_BeatFifoId <= _GEN_923;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1c == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_28_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_28_rvalid <= _GEN_220;
      end
    end else begin
      readStack_28_rvalid <= _GEN_220;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1c == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_28_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1c == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_28_entryid <= _idxInsert_T_62;
        end else begin
          readStack_28_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1c == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_28_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1c == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_28_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1c == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_28_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1c == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_28_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_28_readStatus <= _GEN_348;
      end
    end else begin
      readStack_28_readStatus <= _GEN_348;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1c == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_28_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1c == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_28_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_28 & readStack_28_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_28_entryFifoId <= _readStack_28_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_28_entryFifoId <= _GEN_508;
      end
    end else begin
      readStack_28_entryFifoId <= _GEN_508;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_28_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_28_rvalid & readStack_28_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_28_BeatFifoId <= _readStack_28_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_28_BeatFifoId <= _GEN_924;
      end
    end else begin
      readStack_28_BeatFifoId <= _GEN_924;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1d == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_29_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_29_rvalid <= _GEN_221;
      end
    end else begin
      readStack_29_rvalid <= _GEN_221;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1d == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_29_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1d == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_29_entryid <= _idxInsert_T_62;
        end else begin
          readStack_29_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1d == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_29_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1d == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_29_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1d == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_29_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1d == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_29_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_29_readStatus <= _GEN_349;
      end
    end else begin
      readStack_29_readStatus <= _GEN_349;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1d == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_29_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1d == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_29_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_29 & readStack_29_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_29_entryFifoId <= _readStack_29_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_29_entryFifoId <= _GEN_509;
      end
    end else begin
      readStack_29_entryFifoId <= _GEN_509;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_29_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_29_rvalid & readStack_29_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_29_BeatFifoId <= _readStack_29_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_29_BeatFifoId <= _GEN_925;
      end
    end else begin
      readStack_29_BeatFifoId <= _GEN_925;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1e == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_30_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_30_rvalid <= _GEN_222;
      end
    end else begin
      readStack_30_rvalid <= _GEN_222;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1e == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_30_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1e == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_30_entryid <= _idxInsert_T_62;
        end else begin
          readStack_30_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1e == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_30_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1e == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_30_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1e == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_30_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1e == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_30_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_30_readStatus <= _GEN_350;
      end
    end else begin
      readStack_30_readStatus <= _GEN_350;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1e == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_30_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1e == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_30_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_30 & readStack_30_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_30_entryFifoId <= _readStack_30_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_30_entryFifoId <= _GEN_510;
      end
    end else begin
      readStack_30_entryFifoId <= _GEN_510;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_30_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_30_rvalid & readStack_30_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_30_BeatFifoId <= _readStack_30_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_30_BeatFifoId <= _GEN_926;
      end
    end else begin
      readStack_30_BeatFifoId <= _GEN_926;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_rvalid <= 1'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (5'h1f == axirespArb_io_chosen) begin // @[ReadStack.scala 192:36]
        readStack_31_rvalid <= 1'h0; // @[ReadStack.scala 192:36]
      end else begin
        readStack_31_rvalid <= _GEN_223;
      end
    end else begin
      readStack_31_rvalid <= _GEN_223;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_raddress <= 35'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1f == idxInsert) begin // @[ReadStack.scala 85:22]
        readStack_31_raddress <= io_axiReq_in_ar_bits_addr; // @[ReadStack.scala 85:22]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_entryid <= 5'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1f == idxInsert) begin // @[ReadStack.scala 84:21]
        if (alloc) begin // @[ReadStack.scala 74:22]
          readStack_31_entryid <= _idxInsert_T_62;
        end else begin
          readStack_31_entryid <= 5'h0;
        end
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_arid <= 14'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1f == idxInsert) begin // @[ReadStack.scala 86:18]
        readStack_31_arid <= io_axiReq_in_ar_bits_id; // @[ReadStack.scala 86:18]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_ardata <= 256'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1f == respEntryId) begin // @[ReadStack.scala 155:20]
      readStack_31_ardata <= io_tlResp_in_d_bits_data; // @[ReadStack.scala 155:20]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_readStatus <= 2'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1f == respEntryId) begin // @[ReadStack.scala 156:24]
      readStack_31_readStatus <= 2'h3; // @[ReadStack.scala 156:24]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (5'h1f == axireqArb_io_chosen) begin // @[ReadStack.scala 140:34]
        readStack_31_readStatus <= 2'h2; // @[ReadStack.scala 140:34]
      end else begin
        readStack_31_readStatus <= _GEN_351;
      end
    end else begin
      readStack_31_readStatus <= _GEN_351;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_respStatus <= 4'h0; // @[ReadStack.scala 63:26]
    end else if (5'h1f == respEntryId) begin // @[ReadStack.scala 157:24]
      readStack_31_respStatus <= _readStack_respEntryId_respStatus; // @[ReadStack.scala 157:24]
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_rsize <= 8'h0; // @[ReadStack.scala 63:26]
    end else if (alloc) begin // @[ReadStack.scala 78:5]
      if (5'h1f == idxInsert) begin // @[ReadStack.scala 88:19]
        readStack_31_rsize <= r_size1[7:0]; // @[ReadStack.scala 88:19]
      end
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_entryFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_1) begin // @[ReadStack.scala 139:3]
      if (_hasWaitTLReq_T_31 & readStack_31_rvalid) begin // @[ReadStack.scala 143:51]
        readStack_31_entryFifoId <= _readStack_31_entryFifoId_T_1; // @[ReadStack.scala 144:23]
      end else begin
        readStack_31_entryFifoId <= _GEN_511;
      end
    end else begin
      readStack_31_entryFifoId <= _GEN_511;
    end
    if (reset) begin // @[ReadStack.scala 63:26]
      readStack_31_BeatFifoId <= 6'h0; // @[ReadStack.scala 63:26]
    end else if (_T_72) begin // @[ReadStack.scala 191:30]
      if (readStack_31_rvalid & readStack_31_arid == _GEN_1023) begin // @[ReadStack.scala 196:67]
        readStack_31_BeatFifoId <= _readStack_31_BeatFifoId_T_1; // @[ReadStack.scala 197:26]
      end else begin
        readStack_31_BeatFifoId <= _GEN_927;
      end
    end else begin
      readStack_31_BeatFifoId <= _GEN_927;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  readStack_0_rvalid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  readStack_0_raddress = _RAND_1[34:0];
  _RAND_2 = {1{`RANDOM}};
  readStack_0_entryid = _RAND_2[4:0];
  _RAND_3 = {1{`RANDOM}};
  readStack_0_arid = _RAND_3[13:0];
  _RAND_4 = {8{`RANDOM}};
  readStack_0_ardata = _RAND_4[255:0];
  _RAND_5 = {1{`RANDOM}};
  readStack_0_readStatus = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  readStack_0_respStatus = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  readStack_0_rsize = _RAND_7[7:0];
  _RAND_8 = {1{`RANDOM}};
  readStack_0_entryFifoId = _RAND_8[5:0];
  _RAND_9 = {1{`RANDOM}};
  readStack_0_BeatFifoId = _RAND_9[5:0];
  _RAND_10 = {1{`RANDOM}};
  readStack_1_rvalid = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  readStack_1_raddress = _RAND_11[34:0];
  _RAND_12 = {1{`RANDOM}};
  readStack_1_entryid = _RAND_12[4:0];
  _RAND_13 = {1{`RANDOM}};
  readStack_1_arid = _RAND_13[13:0];
  _RAND_14 = {8{`RANDOM}};
  readStack_1_ardata = _RAND_14[255:0];
  _RAND_15 = {1{`RANDOM}};
  readStack_1_readStatus = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  readStack_1_respStatus = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  readStack_1_rsize = _RAND_17[7:0];
  _RAND_18 = {1{`RANDOM}};
  readStack_1_entryFifoId = _RAND_18[5:0];
  _RAND_19 = {1{`RANDOM}};
  readStack_1_BeatFifoId = _RAND_19[5:0];
  _RAND_20 = {1{`RANDOM}};
  readStack_2_rvalid = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  readStack_2_raddress = _RAND_21[34:0];
  _RAND_22 = {1{`RANDOM}};
  readStack_2_entryid = _RAND_22[4:0];
  _RAND_23 = {1{`RANDOM}};
  readStack_2_arid = _RAND_23[13:0];
  _RAND_24 = {8{`RANDOM}};
  readStack_2_ardata = _RAND_24[255:0];
  _RAND_25 = {1{`RANDOM}};
  readStack_2_readStatus = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  readStack_2_respStatus = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  readStack_2_rsize = _RAND_27[7:0];
  _RAND_28 = {1{`RANDOM}};
  readStack_2_entryFifoId = _RAND_28[5:0];
  _RAND_29 = {1{`RANDOM}};
  readStack_2_BeatFifoId = _RAND_29[5:0];
  _RAND_30 = {1{`RANDOM}};
  readStack_3_rvalid = _RAND_30[0:0];
  _RAND_31 = {2{`RANDOM}};
  readStack_3_raddress = _RAND_31[34:0];
  _RAND_32 = {1{`RANDOM}};
  readStack_3_entryid = _RAND_32[4:0];
  _RAND_33 = {1{`RANDOM}};
  readStack_3_arid = _RAND_33[13:0];
  _RAND_34 = {8{`RANDOM}};
  readStack_3_ardata = _RAND_34[255:0];
  _RAND_35 = {1{`RANDOM}};
  readStack_3_readStatus = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  readStack_3_respStatus = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  readStack_3_rsize = _RAND_37[7:0];
  _RAND_38 = {1{`RANDOM}};
  readStack_3_entryFifoId = _RAND_38[5:0];
  _RAND_39 = {1{`RANDOM}};
  readStack_3_BeatFifoId = _RAND_39[5:0];
  _RAND_40 = {1{`RANDOM}};
  readStack_4_rvalid = _RAND_40[0:0];
  _RAND_41 = {2{`RANDOM}};
  readStack_4_raddress = _RAND_41[34:0];
  _RAND_42 = {1{`RANDOM}};
  readStack_4_entryid = _RAND_42[4:0];
  _RAND_43 = {1{`RANDOM}};
  readStack_4_arid = _RAND_43[13:0];
  _RAND_44 = {8{`RANDOM}};
  readStack_4_ardata = _RAND_44[255:0];
  _RAND_45 = {1{`RANDOM}};
  readStack_4_readStatus = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  readStack_4_respStatus = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  readStack_4_rsize = _RAND_47[7:0];
  _RAND_48 = {1{`RANDOM}};
  readStack_4_entryFifoId = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  readStack_4_BeatFifoId = _RAND_49[5:0];
  _RAND_50 = {1{`RANDOM}};
  readStack_5_rvalid = _RAND_50[0:0];
  _RAND_51 = {2{`RANDOM}};
  readStack_5_raddress = _RAND_51[34:0];
  _RAND_52 = {1{`RANDOM}};
  readStack_5_entryid = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  readStack_5_arid = _RAND_53[13:0];
  _RAND_54 = {8{`RANDOM}};
  readStack_5_ardata = _RAND_54[255:0];
  _RAND_55 = {1{`RANDOM}};
  readStack_5_readStatus = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  readStack_5_respStatus = _RAND_56[3:0];
  _RAND_57 = {1{`RANDOM}};
  readStack_5_rsize = _RAND_57[7:0];
  _RAND_58 = {1{`RANDOM}};
  readStack_5_entryFifoId = _RAND_58[5:0];
  _RAND_59 = {1{`RANDOM}};
  readStack_5_BeatFifoId = _RAND_59[5:0];
  _RAND_60 = {1{`RANDOM}};
  readStack_6_rvalid = _RAND_60[0:0];
  _RAND_61 = {2{`RANDOM}};
  readStack_6_raddress = _RAND_61[34:0];
  _RAND_62 = {1{`RANDOM}};
  readStack_6_entryid = _RAND_62[4:0];
  _RAND_63 = {1{`RANDOM}};
  readStack_6_arid = _RAND_63[13:0];
  _RAND_64 = {8{`RANDOM}};
  readStack_6_ardata = _RAND_64[255:0];
  _RAND_65 = {1{`RANDOM}};
  readStack_6_readStatus = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  readStack_6_respStatus = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  readStack_6_rsize = _RAND_67[7:0];
  _RAND_68 = {1{`RANDOM}};
  readStack_6_entryFifoId = _RAND_68[5:0];
  _RAND_69 = {1{`RANDOM}};
  readStack_6_BeatFifoId = _RAND_69[5:0];
  _RAND_70 = {1{`RANDOM}};
  readStack_7_rvalid = _RAND_70[0:0];
  _RAND_71 = {2{`RANDOM}};
  readStack_7_raddress = _RAND_71[34:0];
  _RAND_72 = {1{`RANDOM}};
  readStack_7_entryid = _RAND_72[4:0];
  _RAND_73 = {1{`RANDOM}};
  readStack_7_arid = _RAND_73[13:0];
  _RAND_74 = {8{`RANDOM}};
  readStack_7_ardata = _RAND_74[255:0];
  _RAND_75 = {1{`RANDOM}};
  readStack_7_readStatus = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  readStack_7_respStatus = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  readStack_7_rsize = _RAND_77[7:0];
  _RAND_78 = {1{`RANDOM}};
  readStack_7_entryFifoId = _RAND_78[5:0];
  _RAND_79 = {1{`RANDOM}};
  readStack_7_BeatFifoId = _RAND_79[5:0];
  _RAND_80 = {1{`RANDOM}};
  readStack_8_rvalid = _RAND_80[0:0];
  _RAND_81 = {2{`RANDOM}};
  readStack_8_raddress = _RAND_81[34:0];
  _RAND_82 = {1{`RANDOM}};
  readStack_8_entryid = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  readStack_8_arid = _RAND_83[13:0];
  _RAND_84 = {8{`RANDOM}};
  readStack_8_ardata = _RAND_84[255:0];
  _RAND_85 = {1{`RANDOM}};
  readStack_8_readStatus = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  readStack_8_respStatus = _RAND_86[3:0];
  _RAND_87 = {1{`RANDOM}};
  readStack_8_rsize = _RAND_87[7:0];
  _RAND_88 = {1{`RANDOM}};
  readStack_8_entryFifoId = _RAND_88[5:0];
  _RAND_89 = {1{`RANDOM}};
  readStack_8_BeatFifoId = _RAND_89[5:0];
  _RAND_90 = {1{`RANDOM}};
  readStack_9_rvalid = _RAND_90[0:0];
  _RAND_91 = {2{`RANDOM}};
  readStack_9_raddress = _RAND_91[34:0];
  _RAND_92 = {1{`RANDOM}};
  readStack_9_entryid = _RAND_92[4:0];
  _RAND_93 = {1{`RANDOM}};
  readStack_9_arid = _RAND_93[13:0];
  _RAND_94 = {8{`RANDOM}};
  readStack_9_ardata = _RAND_94[255:0];
  _RAND_95 = {1{`RANDOM}};
  readStack_9_readStatus = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  readStack_9_respStatus = _RAND_96[3:0];
  _RAND_97 = {1{`RANDOM}};
  readStack_9_rsize = _RAND_97[7:0];
  _RAND_98 = {1{`RANDOM}};
  readStack_9_entryFifoId = _RAND_98[5:0];
  _RAND_99 = {1{`RANDOM}};
  readStack_9_BeatFifoId = _RAND_99[5:0];
  _RAND_100 = {1{`RANDOM}};
  readStack_10_rvalid = _RAND_100[0:0];
  _RAND_101 = {2{`RANDOM}};
  readStack_10_raddress = _RAND_101[34:0];
  _RAND_102 = {1{`RANDOM}};
  readStack_10_entryid = _RAND_102[4:0];
  _RAND_103 = {1{`RANDOM}};
  readStack_10_arid = _RAND_103[13:0];
  _RAND_104 = {8{`RANDOM}};
  readStack_10_ardata = _RAND_104[255:0];
  _RAND_105 = {1{`RANDOM}};
  readStack_10_readStatus = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  readStack_10_respStatus = _RAND_106[3:0];
  _RAND_107 = {1{`RANDOM}};
  readStack_10_rsize = _RAND_107[7:0];
  _RAND_108 = {1{`RANDOM}};
  readStack_10_entryFifoId = _RAND_108[5:0];
  _RAND_109 = {1{`RANDOM}};
  readStack_10_BeatFifoId = _RAND_109[5:0];
  _RAND_110 = {1{`RANDOM}};
  readStack_11_rvalid = _RAND_110[0:0];
  _RAND_111 = {2{`RANDOM}};
  readStack_11_raddress = _RAND_111[34:0];
  _RAND_112 = {1{`RANDOM}};
  readStack_11_entryid = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  readStack_11_arid = _RAND_113[13:0];
  _RAND_114 = {8{`RANDOM}};
  readStack_11_ardata = _RAND_114[255:0];
  _RAND_115 = {1{`RANDOM}};
  readStack_11_readStatus = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  readStack_11_respStatus = _RAND_116[3:0];
  _RAND_117 = {1{`RANDOM}};
  readStack_11_rsize = _RAND_117[7:0];
  _RAND_118 = {1{`RANDOM}};
  readStack_11_entryFifoId = _RAND_118[5:0];
  _RAND_119 = {1{`RANDOM}};
  readStack_11_BeatFifoId = _RAND_119[5:0];
  _RAND_120 = {1{`RANDOM}};
  readStack_12_rvalid = _RAND_120[0:0];
  _RAND_121 = {2{`RANDOM}};
  readStack_12_raddress = _RAND_121[34:0];
  _RAND_122 = {1{`RANDOM}};
  readStack_12_entryid = _RAND_122[4:0];
  _RAND_123 = {1{`RANDOM}};
  readStack_12_arid = _RAND_123[13:0];
  _RAND_124 = {8{`RANDOM}};
  readStack_12_ardata = _RAND_124[255:0];
  _RAND_125 = {1{`RANDOM}};
  readStack_12_readStatus = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  readStack_12_respStatus = _RAND_126[3:0];
  _RAND_127 = {1{`RANDOM}};
  readStack_12_rsize = _RAND_127[7:0];
  _RAND_128 = {1{`RANDOM}};
  readStack_12_entryFifoId = _RAND_128[5:0];
  _RAND_129 = {1{`RANDOM}};
  readStack_12_BeatFifoId = _RAND_129[5:0];
  _RAND_130 = {1{`RANDOM}};
  readStack_13_rvalid = _RAND_130[0:0];
  _RAND_131 = {2{`RANDOM}};
  readStack_13_raddress = _RAND_131[34:0];
  _RAND_132 = {1{`RANDOM}};
  readStack_13_entryid = _RAND_132[4:0];
  _RAND_133 = {1{`RANDOM}};
  readStack_13_arid = _RAND_133[13:0];
  _RAND_134 = {8{`RANDOM}};
  readStack_13_ardata = _RAND_134[255:0];
  _RAND_135 = {1{`RANDOM}};
  readStack_13_readStatus = _RAND_135[1:0];
  _RAND_136 = {1{`RANDOM}};
  readStack_13_respStatus = _RAND_136[3:0];
  _RAND_137 = {1{`RANDOM}};
  readStack_13_rsize = _RAND_137[7:0];
  _RAND_138 = {1{`RANDOM}};
  readStack_13_entryFifoId = _RAND_138[5:0];
  _RAND_139 = {1{`RANDOM}};
  readStack_13_BeatFifoId = _RAND_139[5:0];
  _RAND_140 = {1{`RANDOM}};
  readStack_14_rvalid = _RAND_140[0:0];
  _RAND_141 = {2{`RANDOM}};
  readStack_14_raddress = _RAND_141[34:0];
  _RAND_142 = {1{`RANDOM}};
  readStack_14_entryid = _RAND_142[4:0];
  _RAND_143 = {1{`RANDOM}};
  readStack_14_arid = _RAND_143[13:0];
  _RAND_144 = {8{`RANDOM}};
  readStack_14_ardata = _RAND_144[255:0];
  _RAND_145 = {1{`RANDOM}};
  readStack_14_readStatus = _RAND_145[1:0];
  _RAND_146 = {1{`RANDOM}};
  readStack_14_respStatus = _RAND_146[3:0];
  _RAND_147 = {1{`RANDOM}};
  readStack_14_rsize = _RAND_147[7:0];
  _RAND_148 = {1{`RANDOM}};
  readStack_14_entryFifoId = _RAND_148[5:0];
  _RAND_149 = {1{`RANDOM}};
  readStack_14_BeatFifoId = _RAND_149[5:0];
  _RAND_150 = {1{`RANDOM}};
  readStack_15_rvalid = _RAND_150[0:0];
  _RAND_151 = {2{`RANDOM}};
  readStack_15_raddress = _RAND_151[34:0];
  _RAND_152 = {1{`RANDOM}};
  readStack_15_entryid = _RAND_152[4:0];
  _RAND_153 = {1{`RANDOM}};
  readStack_15_arid = _RAND_153[13:0];
  _RAND_154 = {8{`RANDOM}};
  readStack_15_ardata = _RAND_154[255:0];
  _RAND_155 = {1{`RANDOM}};
  readStack_15_readStatus = _RAND_155[1:0];
  _RAND_156 = {1{`RANDOM}};
  readStack_15_respStatus = _RAND_156[3:0];
  _RAND_157 = {1{`RANDOM}};
  readStack_15_rsize = _RAND_157[7:0];
  _RAND_158 = {1{`RANDOM}};
  readStack_15_entryFifoId = _RAND_158[5:0];
  _RAND_159 = {1{`RANDOM}};
  readStack_15_BeatFifoId = _RAND_159[5:0];
  _RAND_160 = {1{`RANDOM}};
  readStack_16_rvalid = _RAND_160[0:0];
  _RAND_161 = {2{`RANDOM}};
  readStack_16_raddress = _RAND_161[34:0];
  _RAND_162 = {1{`RANDOM}};
  readStack_16_entryid = _RAND_162[4:0];
  _RAND_163 = {1{`RANDOM}};
  readStack_16_arid = _RAND_163[13:0];
  _RAND_164 = {8{`RANDOM}};
  readStack_16_ardata = _RAND_164[255:0];
  _RAND_165 = {1{`RANDOM}};
  readStack_16_readStatus = _RAND_165[1:0];
  _RAND_166 = {1{`RANDOM}};
  readStack_16_respStatus = _RAND_166[3:0];
  _RAND_167 = {1{`RANDOM}};
  readStack_16_rsize = _RAND_167[7:0];
  _RAND_168 = {1{`RANDOM}};
  readStack_16_entryFifoId = _RAND_168[5:0];
  _RAND_169 = {1{`RANDOM}};
  readStack_16_BeatFifoId = _RAND_169[5:0];
  _RAND_170 = {1{`RANDOM}};
  readStack_17_rvalid = _RAND_170[0:0];
  _RAND_171 = {2{`RANDOM}};
  readStack_17_raddress = _RAND_171[34:0];
  _RAND_172 = {1{`RANDOM}};
  readStack_17_entryid = _RAND_172[4:0];
  _RAND_173 = {1{`RANDOM}};
  readStack_17_arid = _RAND_173[13:0];
  _RAND_174 = {8{`RANDOM}};
  readStack_17_ardata = _RAND_174[255:0];
  _RAND_175 = {1{`RANDOM}};
  readStack_17_readStatus = _RAND_175[1:0];
  _RAND_176 = {1{`RANDOM}};
  readStack_17_respStatus = _RAND_176[3:0];
  _RAND_177 = {1{`RANDOM}};
  readStack_17_rsize = _RAND_177[7:0];
  _RAND_178 = {1{`RANDOM}};
  readStack_17_entryFifoId = _RAND_178[5:0];
  _RAND_179 = {1{`RANDOM}};
  readStack_17_BeatFifoId = _RAND_179[5:0];
  _RAND_180 = {1{`RANDOM}};
  readStack_18_rvalid = _RAND_180[0:0];
  _RAND_181 = {2{`RANDOM}};
  readStack_18_raddress = _RAND_181[34:0];
  _RAND_182 = {1{`RANDOM}};
  readStack_18_entryid = _RAND_182[4:0];
  _RAND_183 = {1{`RANDOM}};
  readStack_18_arid = _RAND_183[13:0];
  _RAND_184 = {8{`RANDOM}};
  readStack_18_ardata = _RAND_184[255:0];
  _RAND_185 = {1{`RANDOM}};
  readStack_18_readStatus = _RAND_185[1:0];
  _RAND_186 = {1{`RANDOM}};
  readStack_18_respStatus = _RAND_186[3:0];
  _RAND_187 = {1{`RANDOM}};
  readStack_18_rsize = _RAND_187[7:0];
  _RAND_188 = {1{`RANDOM}};
  readStack_18_entryFifoId = _RAND_188[5:0];
  _RAND_189 = {1{`RANDOM}};
  readStack_18_BeatFifoId = _RAND_189[5:0];
  _RAND_190 = {1{`RANDOM}};
  readStack_19_rvalid = _RAND_190[0:0];
  _RAND_191 = {2{`RANDOM}};
  readStack_19_raddress = _RAND_191[34:0];
  _RAND_192 = {1{`RANDOM}};
  readStack_19_entryid = _RAND_192[4:0];
  _RAND_193 = {1{`RANDOM}};
  readStack_19_arid = _RAND_193[13:0];
  _RAND_194 = {8{`RANDOM}};
  readStack_19_ardata = _RAND_194[255:0];
  _RAND_195 = {1{`RANDOM}};
  readStack_19_readStatus = _RAND_195[1:0];
  _RAND_196 = {1{`RANDOM}};
  readStack_19_respStatus = _RAND_196[3:0];
  _RAND_197 = {1{`RANDOM}};
  readStack_19_rsize = _RAND_197[7:0];
  _RAND_198 = {1{`RANDOM}};
  readStack_19_entryFifoId = _RAND_198[5:0];
  _RAND_199 = {1{`RANDOM}};
  readStack_19_BeatFifoId = _RAND_199[5:0];
  _RAND_200 = {1{`RANDOM}};
  readStack_20_rvalid = _RAND_200[0:0];
  _RAND_201 = {2{`RANDOM}};
  readStack_20_raddress = _RAND_201[34:0];
  _RAND_202 = {1{`RANDOM}};
  readStack_20_entryid = _RAND_202[4:0];
  _RAND_203 = {1{`RANDOM}};
  readStack_20_arid = _RAND_203[13:0];
  _RAND_204 = {8{`RANDOM}};
  readStack_20_ardata = _RAND_204[255:0];
  _RAND_205 = {1{`RANDOM}};
  readStack_20_readStatus = _RAND_205[1:0];
  _RAND_206 = {1{`RANDOM}};
  readStack_20_respStatus = _RAND_206[3:0];
  _RAND_207 = {1{`RANDOM}};
  readStack_20_rsize = _RAND_207[7:0];
  _RAND_208 = {1{`RANDOM}};
  readStack_20_entryFifoId = _RAND_208[5:0];
  _RAND_209 = {1{`RANDOM}};
  readStack_20_BeatFifoId = _RAND_209[5:0];
  _RAND_210 = {1{`RANDOM}};
  readStack_21_rvalid = _RAND_210[0:0];
  _RAND_211 = {2{`RANDOM}};
  readStack_21_raddress = _RAND_211[34:0];
  _RAND_212 = {1{`RANDOM}};
  readStack_21_entryid = _RAND_212[4:0];
  _RAND_213 = {1{`RANDOM}};
  readStack_21_arid = _RAND_213[13:0];
  _RAND_214 = {8{`RANDOM}};
  readStack_21_ardata = _RAND_214[255:0];
  _RAND_215 = {1{`RANDOM}};
  readStack_21_readStatus = _RAND_215[1:0];
  _RAND_216 = {1{`RANDOM}};
  readStack_21_respStatus = _RAND_216[3:0];
  _RAND_217 = {1{`RANDOM}};
  readStack_21_rsize = _RAND_217[7:0];
  _RAND_218 = {1{`RANDOM}};
  readStack_21_entryFifoId = _RAND_218[5:0];
  _RAND_219 = {1{`RANDOM}};
  readStack_21_BeatFifoId = _RAND_219[5:0];
  _RAND_220 = {1{`RANDOM}};
  readStack_22_rvalid = _RAND_220[0:0];
  _RAND_221 = {2{`RANDOM}};
  readStack_22_raddress = _RAND_221[34:0];
  _RAND_222 = {1{`RANDOM}};
  readStack_22_entryid = _RAND_222[4:0];
  _RAND_223 = {1{`RANDOM}};
  readStack_22_arid = _RAND_223[13:0];
  _RAND_224 = {8{`RANDOM}};
  readStack_22_ardata = _RAND_224[255:0];
  _RAND_225 = {1{`RANDOM}};
  readStack_22_readStatus = _RAND_225[1:0];
  _RAND_226 = {1{`RANDOM}};
  readStack_22_respStatus = _RAND_226[3:0];
  _RAND_227 = {1{`RANDOM}};
  readStack_22_rsize = _RAND_227[7:0];
  _RAND_228 = {1{`RANDOM}};
  readStack_22_entryFifoId = _RAND_228[5:0];
  _RAND_229 = {1{`RANDOM}};
  readStack_22_BeatFifoId = _RAND_229[5:0];
  _RAND_230 = {1{`RANDOM}};
  readStack_23_rvalid = _RAND_230[0:0];
  _RAND_231 = {2{`RANDOM}};
  readStack_23_raddress = _RAND_231[34:0];
  _RAND_232 = {1{`RANDOM}};
  readStack_23_entryid = _RAND_232[4:0];
  _RAND_233 = {1{`RANDOM}};
  readStack_23_arid = _RAND_233[13:0];
  _RAND_234 = {8{`RANDOM}};
  readStack_23_ardata = _RAND_234[255:0];
  _RAND_235 = {1{`RANDOM}};
  readStack_23_readStatus = _RAND_235[1:0];
  _RAND_236 = {1{`RANDOM}};
  readStack_23_respStatus = _RAND_236[3:0];
  _RAND_237 = {1{`RANDOM}};
  readStack_23_rsize = _RAND_237[7:0];
  _RAND_238 = {1{`RANDOM}};
  readStack_23_entryFifoId = _RAND_238[5:0];
  _RAND_239 = {1{`RANDOM}};
  readStack_23_BeatFifoId = _RAND_239[5:0];
  _RAND_240 = {1{`RANDOM}};
  readStack_24_rvalid = _RAND_240[0:0];
  _RAND_241 = {2{`RANDOM}};
  readStack_24_raddress = _RAND_241[34:0];
  _RAND_242 = {1{`RANDOM}};
  readStack_24_entryid = _RAND_242[4:0];
  _RAND_243 = {1{`RANDOM}};
  readStack_24_arid = _RAND_243[13:0];
  _RAND_244 = {8{`RANDOM}};
  readStack_24_ardata = _RAND_244[255:0];
  _RAND_245 = {1{`RANDOM}};
  readStack_24_readStatus = _RAND_245[1:0];
  _RAND_246 = {1{`RANDOM}};
  readStack_24_respStatus = _RAND_246[3:0];
  _RAND_247 = {1{`RANDOM}};
  readStack_24_rsize = _RAND_247[7:0];
  _RAND_248 = {1{`RANDOM}};
  readStack_24_entryFifoId = _RAND_248[5:0];
  _RAND_249 = {1{`RANDOM}};
  readStack_24_BeatFifoId = _RAND_249[5:0];
  _RAND_250 = {1{`RANDOM}};
  readStack_25_rvalid = _RAND_250[0:0];
  _RAND_251 = {2{`RANDOM}};
  readStack_25_raddress = _RAND_251[34:0];
  _RAND_252 = {1{`RANDOM}};
  readStack_25_entryid = _RAND_252[4:0];
  _RAND_253 = {1{`RANDOM}};
  readStack_25_arid = _RAND_253[13:0];
  _RAND_254 = {8{`RANDOM}};
  readStack_25_ardata = _RAND_254[255:0];
  _RAND_255 = {1{`RANDOM}};
  readStack_25_readStatus = _RAND_255[1:0];
  _RAND_256 = {1{`RANDOM}};
  readStack_25_respStatus = _RAND_256[3:0];
  _RAND_257 = {1{`RANDOM}};
  readStack_25_rsize = _RAND_257[7:0];
  _RAND_258 = {1{`RANDOM}};
  readStack_25_entryFifoId = _RAND_258[5:0];
  _RAND_259 = {1{`RANDOM}};
  readStack_25_BeatFifoId = _RAND_259[5:0];
  _RAND_260 = {1{`RANDOM}};
  readStack_26_rvalid = _RAND_260[0:0];
  _RAND_261 = {2{`RANDOM}};
  readStack_26_raddress = _RAND_261[34:0];
  _RAND_262 = {1{`RANDOM}};
  readStack_26_entryid = _RAND_262[4:0];
  _RAND_263 = {1{`RANDOM}};
  readStack_26_arid = _RAND_263[13:0];
  _RAND_264 = {8{`RANDOM}};
  readStack_26_ardata = _RAND_264[255:0];
  _RAND_265 = {1{`RANDOM}};
  readStack_26_readStatus = _RAND_265[1:0];
  _RAND_266 = {1{`RANDOM}};
  readStack_26_respStatus = _RAND_266[3:0];
  _RAND_267 = {1{`RANDOM}};
  readStack_26_rsize = _RAND_267[7:0];
  _RAND_268 = {1{`RANDOM}};
  readStack_26_entryFifoId = _RAND_268[5:0];
  _RAND_269 = {1{`RANDOM}};
  readStack_26_BeatFifoId = _RAND_269[5:0];
  _RAND_270 = {1{`RANDOM}};
  readStack_27_rvalid = _RAND_270[0:0];
  _RAND_271 = {2{`RANDOM}};
  readStack_27_raddress = _RAND_271[34:0];
  _RAND_272 = {1{`RANDOM}};
  readStack_27_entryid = _RAND_272[4:0];
  _RAND_273 = {1{`RANDOM}};
  readStack_27_arid = _RAND_273[13:0];
  _RAND_274 = {8{`RANDOM}};
  readStack_27_ardata = _RAND_274[255:0];
  _RAND_275 = {1{`RANDOM}};
  readStack_27_readStatus = _RAND_275[1:0];
  _RAND_276 = {1{`RANDOM}};
  readStack_27_respStatus = _RAND_276[3:0];
  _RAND_277 = {1{`RANDOM}};
  readStack_27_rsize = _RAND_277[7:0];
  _RAND_278 = {1{`RANDOM}};
  readStack_27_entryFifoId = _RAND_278[5:0];
  _RAND_279 = {1{`RANDOM}};
  readStack_27_BeatFifoId = _RAND_279[5:0];
  _RAND_280 = {1{`RANDOM}};
  readStack_28_rvalid = _RAND_280[0:0];
  _RAND_281 = {2{`RANDOM}};
  readStack_28_raddress = _RAND_281[34:0];
  _RAND_282 = {1{`RANDOM}};
  readStack_28_entryid = _RAND_282[4:0];
  _RAND_283 = {1{`RANDOM}};
  readStack_28_arid = _RAND_283[13:0];
  _RAND_284 = {8{`RANDOM}};
  readStack_28_ardata = _RAND_284[255:0];
  _RAND_285 = {1{`RANDOM}};
  readStack_28_readStatus = _RAND_285[1:0];
  _RAND_286 = {1{`RANDOM}};
  readStack_28_respStatus = _RAND_286[3:0];
  _RAND_287 = {1{`RANDOM}};
  readStack_28_rsize = _RAND_287[7:0];
  _RAND_288 = {1{`RANDOM}};
  readStack_28_entryFifoId = _RAND_288[5:0];
  _RAND_289 = {1{`RANDOM}};
  readStack_28_BeatFifoId = _RAND_289[5:0];
  _RAND_290 = {1{`RANDOM}};
  readStack_29_rvalid = _RAND_290[0:0];
  _RAND_291 = {2{`RANDOM}};
  readStack_29_raddress = _RAND_291[34:0];
  _RAND_292 = {1{`RANDOM}};
  readStack_29_entryid = _RAND_292[4:0];
  _RAND_293 = {1{`RANDOM}};
  readStack_29_arid = _RAND_293[13:0];
  _RAND_294 = {8{`RANDOM}};
  readStack_29_ardata = _RAND_294[255:0];
  _RAND_295 = {1{`RANDOM}};
  readStack_29_readStatus = _RAND_295[1:0];
  _RAND_296 = {1{`RANDOM}};
  readStack_29_respStatus = _RAND_296[3:0];
  _RAND_297 = {1{`RANDOM}};
  readStack_29_rsize = _RAND_297[7:0];
  _RAND_298 = {1{`RANDOM}};
  readStack_29_entryFifoId = _RAND_298[5:0];
  _RAND_299 = {1{`RANDOM}};
  readStack_29_BeatFifoId = _RAND_299[5:0];
  _RAND_300 = {1{`RANDOM}};
  readStack_30_rvalid = _RAND_300[0:0];
  _RAND_301 = {2{`RANDOM}};
  readStack_30_raddress = _RAND_301[34:0];
  _RAND_302 = {1{`RANDOM}};
  readStack_30_entryid = _RAND_302[4:0];
  _RAND_303 = {1{`RANDOM}};
  readStack_30_arid = _RAND_303[13:0];
  _RAND_304 = {8{`RANDOM}};
  readStack_30_ardata = _RAND_304[255:0];
  _RAND_305 = {1{`RANDOM}};
  readStack_30_readStatus = _RAND_305[1:0];
  _RAND_306 = {1{`RANDOM}};
  readStack_30_respStatus = _RAND_306[3:0];
  _RAND_307 = {1{`RANDOM}};
  readStack_30_rsize = _RAND_307[7:0];
  _RAND_308 = {1{`RANDOM}};
  readStack_30_entryFifoId = _RAND_308[5:0];
  _RAND_309 = {1{`RANDOM}};
  readStack_30_BeatFifoId = _RAND_309[5:0];
  _RAND_310 = {1{`RANDOM}};
  readStack_31_rvalid = _RAND_310[0:0];
  _RAND_311 = {2{`RANDOM}};
  readStack_31_raddress = _RAND_311[34:0];
  _RAND_312 = {1{`RANDOM}};
  readStack_31_entryid = _RAND_312[4:0];
  _RAND_313 = {1{`RANDOM}};
  readStack_31_arid = _RAND_313[13:0];
  _RAND_314 = {8{`RANDOM}};
  readStack_31_ardata = _RAND_314[255:0];
  _RAND_315 = {1{`RANDOM}};
  readStack_31_readStatus = _RAND_315[1:0];
  _RAND_316 = {1{`RANDOM}};
  readStack_31_respStatus = _RAND_316[3:0];
  _RAND_317 = {1{`RANDOM}};
  readStack_31_rsize = _RAND_317[7:0];
  _RAND_318 = {1{`RANDOM}};
  readStack_31_entryFifoId = _RAND_318[5:0];
  _RAND_319 = {1{`RANDOM}};
  readStack_31_BeatFifoId = _RAND_319[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
